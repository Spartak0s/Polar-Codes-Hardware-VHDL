library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

entity synt2 is
port( 
	  address1	: in signed (5 downto 0);
	  stoixeio1	: out signed (80-1 downto 0)
);
end synt2;


architecture struct of synt2 is

    type rom_type is array (35 downto 0) of signed (79 downto 0);
    constant stoixeia : rom_type :=("11111111111111111110010011101001100000010011100001111000000000000000000000000000",
"11111111111111111110010001111010011111001001110111100000000000000000000000000000",
"11111111111111111110010000000110000001111000000100000000000000000000000000000000",
"11111111111111111110001110001011100010101110001100100000000000000000000000000000",
"11111111111111111110001100001010100100010101001101111000000000000000000000000000",
"11111111111111111110001010000010100000111101001101100000000000000000000000000000",
"11111111111111111110000111110010100110010000111100110000000000000000000000000000",
"11111111111111111110000101011010001110100000100000111000000000000000000000000000",
"11111111111111111110000010111000010110100100111100000000000000000000000000000000",
"11111111111111111110000000001100000111111100100011110000000000000000000000000000",
"11111111111111111101111101010100001010100010001111000000000000000000000000000000",
"11111111111111111101111010001111010010110110001000000000000000000000000000000000",
"11111111111111111101110110111011110011110100111010001000000000000000000000000000",
"11111111111111111101110011010111110011110101111101010000000000000000000000000000",
"11111111111111111101101111100001000100010010011101110000000000000000000000000000",
"11111111111111111101101011010100111001001100100101000000000000000000000000000000",
"11111111111111111101100110101111111000011101101001111000000000000000000000000000",
"11111111111111111101100001101110000110011011100100010000000000000000000000000000",
"11111111111111111101011100001010010111101111111010010000000000000000000000000000",
"11111111111111111101010101111110010001011000000001000000000000000000000000000000",
"11111111111111111101001111000001101011001101111000011000000000000000000000000000",
"11111111111111111101000111001001101101000001001110011000000000000000000000000000",
"11111111111111111100111110000111111100000010001111101000000000000000000000000000",
"11111111111111111100110011101000001100011010110100100000000000000000000000000000",
"11111111111111111100100111001110001010001110110101100000000000000000000000000000",
"11111111111111111100011000001111010111100100000111011000000000000000000000000000",
"11111111111111111100000101101001101100010111010010000000000000000000000000000000",
"11111111111111111011101101101110110001011011000001111000000000000000000000000000",
"11111111111111111011001101010100010010111011000110110000000000000000000000000000",
"11111111111111111010011101110011100111110011010000010000000000000000000000000000",
"11111111111111111001001110000110010111010111110010110000000000000000000000000000",
"11111111111111110110011001100101001010101001001101110000000000000000000000000000",
"11111111111111101111001011100000001101001100010010010000000000000000000000000000",
"00000000000100010111101101001010001000110011100111000000111011000000000000000000",
"00000000000010001001101000000001001001011001100111101101011111001000000000000000",
"00000000001010111110001110001110111100110100110101101010000101100000000000000000");

begin

stoixeio1<=stoixeia(to_integer((unsigned(address1))));
end struct;

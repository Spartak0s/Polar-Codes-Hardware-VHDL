----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:10:49 02/17/2016 
-- Design Name: 
-- Module Name:    PartialSumGenerator - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.MyPackage.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PartialSumGenerator is
	Port (estimated : in std_logic_vector(N-2 downto 0);
			partial_sums : out s_2d);
end PartialSumGenerator;

architecture Behavioral of PartialSumGenerator is
	--gnal temp : s_2d;
begin
partial_sums(1)(0) <= estimated(0);
partial_sums(1)(1) <= estimated(256);
partial_sums(1)(2) <= estimated(128);
partial_sums(1)(3) <= estimated(384);
partial_sums(1)(4) <= estimated(64);
partial_sums(1)(5) <= estimated(320);
partial_sums(1)(6) <= estimated(192);
partial_sums(1)(7) <= estimated(448);
partial_sums(1)(8) <= estimated(32);
partial_sums(1)(9) <= estimated(288);
partial_sums(1)(10) <= estimated(160);
partial_sums(1)(11) <= estimated(416);
partial_sums(1)(12) <= estimated(96);
partial_sums(1)(13) <= estimated(352);
partial_sums(1)(14) <= estimated(224);
partial_sums(1)(15) <= estimated(480);
partial_sums(1)(16) <= estimated(16);
partial_sums(1)(17) <= estimated(272);
partial_sums(1)(18) <= estimated(144);
partial_sums(1)(19) <= estimated(400);
partial_sums(1)(20) <= estimated(80);
partial_sums(1)(21) <= estimated(336);
partial_sums(1)(22) <= estimated(208);
partial_sums(1)(23) <= estimated(464);
partial_sums(1)(24) <= estimated(48);
partial_sums(1)(25) <= estimated(304);
partial_sums(1)(26) <= estimated(176);
partial_sums(1)(27) <= estimated(432);
partial_sums(1)(28) <= estimated(112);
partial_sums(1)(29) <= estimated(368);
partial_sums(1)(30) <= estimated(240);
partial_sums(1)(31) <= estimated(496);
partial_sums(1)(32) <= estimated(8);
partial_sums(1)(33) <= estimated(264);
partial_sums(1)(34) <= estimated(136);
partial_sums(1)(35) <= estimated(392);
partial_sums(1)(36) <= estimated(72);
partial_sums(1)(37) <= estimated(328);
partial_sums(1)(38) <= estimated(200);
partial_sums(1)(39) <= estimated(456);
partial_sums(1)(40) <= estimated(40);
partial_sums(1)(41) <= estimated(296);
partial_sums(1)(42) <= estimated(168);
partial_sums(1)(43) <= estimated(424);
partial_sums(1)(44) <= estimated(104);
partial_sums(1)(45) <= estimated(360);
partial_sums(1)(46) <= estimated(232);
partial_sums(1)(47) <= estimated(488);
partial_sums(1)(48) <= estimated(24);
partial_sums(1)(49) <= estimated(280);
partial_sums(1)(50) <= estimated(152);
partial_sums(1)(51) <= estimated(408);
partial_sums(1)(52) <= estimated(88);
partial_sums(1)(53) <= estimated(344);
partial_sums(1)(54) <= estimated(216);
partial_sums(1)(55) <= estimated(472);
partial_sums(1)(56) <= estimated(56);
partial_sums(1)(57) <= estimated(312);
partial_sums(1)(58) <= estimated(184);
partial_sums(1)(59) <= estimated(440);
partial_sums(1)(60) <= estimated(120);
partial_sums(1)(61) <= estimated(376);
partial_sums(1)(62) <= estimated(248);
partial_sums(1)(63) <= estimated(504);
partial_sums(1)(64) <= estimated(4);
partial_sums(1)(65) <= estimated(260);
partial_sums(1)(66) <= estimated(132);
partial_sums(1)(67) <= estimated(388);
partial_sums(1)(68) <= estimated(68);
partial_sums(1)(69) <= estimated(324);
partial_sums(1)(70) <= estimated(196);
partial_sums(1)(71) <= estimated(452);
partial_sums(1)(72) <= estimated(36);
partial_sums(1)(73) <= estimated(292);
partial_sums(1)(74) <= estimated(164);
partial_sums(1)(75) <= estimated(420);
partial_sums(1)(76) <= estimated(100);
partial_sums(1)(77) <= estimated(356);
partial_sums(1)(78) <= estimated(228);
partial_sums(1)(79) <= estimated(484);
partial_sums(1)(80) <= estimated(20);
partial_sums(1)(81) <= estimated(276);
partial_sums(1)(82) <= estimated(148);
partial_sums(1)(83) <= estimated(404);
partial_sums(1)(84) <= estimated(84);
partial_sums(1)(85) <= estimated(340);
partial_sums(1)(86) <= estimated(212);
partial_sums(1)(87) <= estimated(468);
partial_sums(1)(88) <= estimated(52);
partial_sums(1)(89) <= estimated(308);
partial_sums(1)(90) <= estimated(180);
partial_sums(1)(91) <= estimated(436);
partial_sums(1)(92) <= estimated(116);
partial_sums(1)(93) <= estimated(372);
partial_sums(1)(94) <= estimated(244);
partial_sums(1)(95) <= estimated(500);
partial_sums(1)(96) <= estimated(12);
partial_sums(1)(97) <= estimated(268);
partial_sums(1)(98) <= estimated(140);
partial_sums(1)(99) <= estimated(396);
partial_sums(1)(100) <= estimated(76);
partial_sums(1)(101) <= estimated(332);
partial_sums(1)(102) <= estimated(204);
partial_sums(1)(103) <= estimated(460);
partial_sums(1)(104) <= estimated(44);
partial_sums(1)(105) <= estimated(300);
partial_sums(1)(106) <= estimated(172);
partial_sums(1)(107) <= estimated(428);
partial_sums(1)(108) <= estimated(108);
partial_sums(1)(109) <= estimated(364);
partial_sums(1)(110) <= estimated(236);
partial_sums(1)(111) <= estimated(492);
partial_sums(1)(112) <= estimated(28);
partial_sums(1)(113) <= estimated(284);
partial_sums(1)(114) <= estimated(156);
partial_sums(1)(115) <= estimated(412);
partial_sums(1)(116) <= estimated(92);
partial_sums(1)(117) <= estimated(348);
partial_sums(1)(118) <= estimated(220);
partial_sums(1)(119) <= estimated(476);
partial_sums(1)(120) <= estimated(60);
partial_sums(1)(121) <= estimated(316);
partial_sums(1)(122) <= estimated(188);
partial_sums(1)(123) <= estimated(444);
partial_sums(1)(124) <= estimated(124);
partial_sums(1)(125) <= estimated(380);
partial_sums(1)(126) <= estimated(252);
partial_sums(1)(127) <= estimated(508);
partial_sums(1)(128) <= estimated(2);
partial_sums(1)(129) <= estimated(258);
partial_sums(1)(130) <= estimated(130);
partial_sums(1)(131) <= estimated(386);
partial_sums(1)(132) <= estimated(66);
partial_sums(1)(133) <= estimated(322);
partial_sums(1)(134) <= estimated(194);
partial_sums(1)(135) <= estimated(450);
partial_sums(1)(136) <= estimated(34);
partial_sums(1)(137) <= estimated(290);
partial_sums(1)(138) <= estimated(162);
partial_sums(1)(139) <= estimated(418);
partial_sums(1)(140) <= estimated(98);
partial_sums(1)(141) <= estimated(354);
partial_sums(1)(142) <= estimated(226);
partial_sums(1)(143) <= estimated(482);
partial_sums(1)(144) <= estimated(18);
partial_sums(1)(145) <= estimated(274);
partial_sums(1)(146) <= estimated(146);
partial_sums(1)(147) <= estimated(402);
partial_sums(1)(148) <= estimated(82);
partial_sums(1)(149) <= estimated(338);
partial_sums(1)(150) <= estimated(210);
partial_sums(1)(151) <= estimated(466);
partial_sums(1)(152) <= estimated(50);
partial_sums(1)(153) <= estimated(306);
partial_sums(1)(154) <= estimated(178);
partial_sums(1)(155) <= estimated(434);
partial_sums(1)(156) <= estimated(114);
partial_sums(1)(157) <= estimated(370);
partial_sums(1)(158) <= estimated(242);
partial_sums(1)(159) <= estimated(498);
partial_sums(1)(160) <= estimated(10);
partial_sums(1)(161) <= estimated(266);
partial_sums(1)(162) <= estimated(138);
partial_sums(1)(163) <= estimated(394);
partial_sums(1)(164) <= estimated(74);
partial_sums(1)(165) <= estimated(330);
partial_sums(1)(166) <= estimated(202);
partial_sums(1)(167) <= estimated(458);
partial_sums(1)(168) <= estimated(42);
partial_sums(1)(169) <= estimated(298);
partial_sums(1)(170) <= estimated(170);
partial_sums(1)(171) <= estimated(426);
partial_sums(1)(172) <= estimated(106);
partial_sums(1)(173) <= estimated(362);
partial_sums(1)(174) <= estimated(234);
partial_sums(1)(175) <= estimated(490);
partial_sums(1)(176) <= estimated(26);
partial_sums(1)(177) <= estimated(282);
partial_sums(1)(178) <= estimated(154);
partial_sums(1)(179) <= estimated(410);
partial_sums(1)(180) <= estimated(90);
partial_sums(1)(181) <= estimated(346);
partial_sums(1)(182) <= estimated(218);
partial_sums(1)(183) <= estimated(474);
partial_sums(1)(184) <= estimated(58);
partial_sums(1)(185) <= estimated(314);
partial_sums(1)(186) <= estimated(186);
partial_sums(1)(187) <= estimated(442);
partial_sums(1)(188) <= estimated(122);
partial_sums(1)(189) <= estimated(378);
partial_sums(1)(190) <= estimated(250);
partial_sums(1)(191) <= estimated(506);
partial_sums(1)(192) <= estimated(6);
partial_sums(1)(193) <= estimated(262);
partial_sums(1)(194) <= estimated(134);
partial_sums(1)(195) <= estimated(390);
partial_sums(1)(196) <= estimated(70);
partial_sums(1)(197) <= estimated(326);
partial_sums(1)(198) <= estimated(198);
partial_sums(1)(199) <= estimated(454);
partial_sums(1)(200) <= estimated(38);
partial_sums(1)(201) <= estimated(294);
partial_sums(1)(202) <= estimated(166);
partial_sums(1)(203) <= estimated(422);
partial_sums(1)(204) <= estimated(102);
partial_sums(1)(205) <= estimated(358);
partial_sums(1)(206) <= estimated(230);
partial_sums(1)(207) <= estimated(486);
partial_sums(1)(208) <= estimated(22);
partial_sums(1)(209) <= estimated(278);
partial_sums(1)(210) <= estimated(150);
partial_sums(1)(211) <= estimated(406);
partial_sums(1)(212) <= estimated(86);
partial_sums(1)(213) <= estimated(342);
partial_sums(1)(214) <= estimated(214);
partial_sums(1)(215) <= estimated(470);
partial_sums(1)(216) <= estimated(54);
partial_sums(1)(217) <= estimated(310);
partial_sums(1)(218) <= estimated(182);
partial_sums(1)(219) <= estimated(438);
partial_sums(1)(220) <= estimated(118);
partial_sums(1)(221) <= estimated(374);
partial_sums(1)(222) <= estimated(246);
partial_sums(1)(223) <= estimated(502);
partial_sums(1)(224) <= estimated(14);
partial_sums(1)(225) <= estimated(270);
partial_sums(1)(226) <= estimated(142);
partial_sums(1)(227) <= estimated(398);
partial_sums(1)(228) <= estimated(78);
partial_sums(1)(229) <= estimated(334);
partial_sums(1)(230) <= estimated(206);
partial_sums(1)(231) <= estimated(462);
partial_sums(1)(232) <= estimated(46);
partial_sums(1)(233) <= estimated(302);
partial_sums(1)(234) <= estimated(174);
partial_sums(1)(235) <= estimated(430);
partial_sums(1)(236) <= estimated(110);
partial_sums(1)(237) <= estimated(366);
partial_sums(1)(238) <= estimated(238);
partial_sums(1)(239) <= estimated(494);
partial_sums(1)(240) <= estimated(30);
partial_sums(1)(241) <= estimated(286);
partial_sums(1)(242) <= estimated(158);
partial_sums(1)(243) <= estimated(414);
partial_sums(1)(244) <= estimated(94);
partial_sums(1)(245) <= estimated(350);
partial_sums(1)(246) <= estimated(222);
partial_sums(1)(247) <= estimated(478);
partial_sums(1)(248) <= estimated(62);
partial_sums(1)(249) <= estimated(318);
partial_sums(1)(250) <= estimated(190);
partial_sums(1)(251) <= estimated(446);
partial_sums(1)(252) <= estimated(126);
partial_sums(1)(253) <= estimated(382);
partial_sums(1)(254) <= estimated(254);
partial_sums(1)(255) <= estimated(510);
partial_sums(2)(0) <= estimated(0) xor estimated(1);
partial_sums(2)(1) <= estimated(256) xor estimated(257);
partial_sums(2)(2) <= estimated(128) xor estimated(129);
partial_sums(2)(3) <= estimated(384) xor estimated(385);
partial_sums(2)(4) <= estimated(64) xor estimated(65);
partial_sums(2)(5) <= estimated(320) xor estimated(321);
partial_sums(2)(6) <= estimated(192) xor estimated(193);
partial_sums(2)(7) <= estimated(448) xor estimated(449);
partial_sums(2)(8) <= estimated(32) xor estimated(33);
partial_sums(2)(9) <= estimated(288) xor estimated(289);
partial_sums(2)(10) <= estimated(160) xor estimated(161);
partial_sums(2)(11) <= estimated(416) xor estimated(417);
partial_sums(2)(12) <= estimated(96) xor estimated(97);
partial_sums(2)(13) <= estimated(352) xor estimated(353);
partial_sums(2)(14) <= estimated(224) xor estimated(225);
partial_sums(2)(15) <= estimated(480) xor estimated(481);
partial_sums(2)(16) <= estimated(16) xor estimated(17);
partial_sums(2)(17) <= estimated(272) xor estimated(273);
partial_sums(2)(18) <= estimated(144) xor estimated(145);
partial_sums(2)(19) <= estimated(400) xor estimated(401);
partial_sums(2)(20) <= estimated(80) xor estimated(81);
partial_sums(2)(21) <= estimated(336) xor estimated(337);
partial_sums(2)(22) <= estimated(208) xor estimated(209);
partial_sums(2)(23) <= estimated(464) xor estimated(465);
partial_sums(2)(24) <= estimated(48) xor estimated(49);
partial_sums(2)(25) <= estimated(304) xor estimated(305);
partial_sums(2)(26) <= estimated(176) xor estimated(177);
partial_sums(2)(27) <= estimated(432) xor estimated(433);
partial_sums(2)(28) <= estimated(112) xor estimated(113);
partial_sums(2)(29) <= estimated(368) xor estimated(369);
partial_sums(2)(30) <= estimated(240) xor estimated(241);
partial_sums(2)(31) <= estimated(496) xor estimated(497);
partial_sums(2)(32) <= estimated(8) xor estimated(9);
partial_sums(2)(33) <= estimated(264) xor estimated(265);
partial_sums(2)(34) <= estimated(136) xor estimated(137);
partial_sums(2)(35) <= estimated(392) xor estimated(393);
partial_sums(2)(36) <= estimated(72) xor estimated(73);
partial_sums(2)(37) <= estimated(328) xor estimated(329);
partial_sums(2)(38) <= estimated(200) xor estimated(201);
partial_sums(2)(39) <= estimated(456) xor estimated(457);
partial_sums(2)(40) <= estimated(40) xor estimated(41);
partial_sums(2)(41) <= estimated(296) xor estimated(297);
partial_sums(2)(42) <= estimated(168) xor estimated(169);
partial_sums(2)(43) <= estimated(424) xor estimated(425);
partial_sums(2)(44) <= estimated(104) xor estimated(105);
partial_sums(2)(45) <= estimated(360) xor estimated(361);
partial_sums(2)(46) <= estimated(232) xor estimated(233);
partial_sums(2)(47) <= estimated(488) xor estimated(489);
partial_sums(2)(48) <= estimated(24) xor estimated(25);
partial_sums(2)(49) <= estimated(280) xor estimated(281);
partial_sums(2)(50) <= estimated(152) xor estimated(153);
partial_sums(2)(51) <= estimated(408) xor estimated(409);
partial_sums(2)(52) <= estimated(88) xor estimated(89);
partial_sums(2)(53) <= estimated(344) xor estimated(345);
partial_sums(2)(54) <= estimated(216) xor estimated(217);
partial_sums(2)(55) <= estimated(472) xor estimated(473);
partial_sums(2)(56) <= estimated(56) xor estimated(57);
partial_sums(2)(57) <= estimated(312) xor estimated(313);
partial_sums(2)(58) <= estimated(184) xor estimated(185);
partial_sums(2)(59) <= estimated(440) xor estimated(441);
partial_sums(2)(60) <= estimated(120) xor estimated(121);
partial_sums(2)(61) <= estimated(376) xor estimated(377);
partial_sums(2)(62) <= estimated(248) xor estimated(249);
partial_sums(2)(63) <= estimated(504) xor estimated(505);
partial_sums(2)(64) <= estimated(4) xor estimated(5);
partial_sums(2)(65) <= estimated(260) xor estimated(261);
partial_sums(2)(66) <= estimated(132) xor estimated(133);
partial_sums(2)(67) <= estimated(388) xor estimated(389);
partial_sums(2)(68) <= estimated(68) xor estimated(69);
partial_sums(2)(69) <= estimated(324) xor estimated(325);
partial_sums(2)(70) <= estimated(196) xor estimated(197);
partial_sums(2)(71) <= estimated(452) xor estimated(453);
partial_sums(2)(72) <= estimated(36) xor estimated(37);
partial_sums(2)(73) <= estimated(292) xor estimated(293);
partial_sums(2)(74) <= estimated(164) xor estimated(165);
partial_sums(2)(75) <= estimated(420) xor estimated(421);
partial_sums(2)(76) <= estimated(100) xor estimated(101);
partial_sums(2)(77) <= estimated(356) xor estimated(357);
partial_sums(2)(78) <= estimated(228) xor estimated(229);
partial_sums(2)(79) <= estimated(484) xor estimated(485);
partial_sums(2)(80) <= estimated(20) xor estimated(21);
partial_sums(2)(81) <= estimated(276) xor estimated(277);
partial_sums(2)(82) <= estimated(148) xor estimated(149);
partial_sums(2)(83) <= estimated(404) xor estimated(405);
partial_sums(2)(84) <= estimated(84) xor estimated(85);
partial_sums(2)(85) <= estimated(340) xor estimated(341);
partial_sums(2)(86) <= estimated(212) xor estimated(213);
partial_sums(2)(87) <= estimated(468) xor estimated(469);
partial_sums(2)(88) <= estimated(52) xor estimated(53);
partial_sums(2)(89) <= estimated(308) xor estimated(309);
partial_sums(2)(90) <= estimated(180) xor estimated(181);
partial_sums(2)(91) <= estimated(436) xor estimated(437);
partial_sums(2)(92) <= estimated(116) xor estimated(117);
partial_sums(2)(93) <= estimated(372) xor estimated(373);
partial_sums(2)(94) <= estimated(244) xor estimated(245);
partial_sums(2)(95) <= estimated(500) xor estimated(501);
partial_sums(2)(96) <= estimated(12) xor estimated(13);
partial_sums(2)(97) <= estimated(268) xor estimated(269);
partial_sums(2)(98) <= estimated(140) xor estimated(141);
partial_sums(2)(99) <= estimated(396) xor estimated(397);
partial_sums(2)(100) <= estimated(76) xor estimated(77);
partial_sums(2)(101) <= estimated(332) xor estimated(333);
partial_sums(2)(102) <= estimated(204) xor estimated(205);
partial_sums(2)(103) <= estimated(460) xor estimated(461);
partial_sums(2)(104) <= estimated(44) xor estimated(45);
partial_sums(2)(105) <= estimated(300) xor estimated(301);
partial_sums(2)(106) <= estimated(172) xor estimated(173);
partial_sums(2)(107) <= estimated(428) xor estimated(429);
partial_sums(2)(108) <= estimated(108) xor estimated(109);
partial_sums(2)(109) <= estimated(364) xor estimated(365);
partial_sums(2)(110) <= estimated(236) xor estimated(237);
partial_sums(2)(111) <= estimated(492) xor estimated(493);
partial_sums(2)(112) <= estimated(28) xor estimated(29);
partial_sums(2)(113) <= estimated(284) xor estimated(285);
partial_sums(2)(114) <= estimated(156) xor estimated(157);
partial_sums(2)(115) <= estimated(412) xor estimated(413);
partial_sums(2)(116) <= estimated(92) xor estimated(93);
partial_sums(2)(117) <= estimated(348) xor estimated(349);
partial_sums(2)(118) <= estimated(220) xor estimated(221);
partial_sums(2)(119) <= estimated(476) xor estimated(477);
partial_sums(2)(120) <= estimated(60) xor estimated(61);
partial_sums(2)(121) <= estimated(316) xor estimated(317);
partial_sums(2)(122) <= estimated(188) xor estimated(189);
partial_sums(2)(123) <= estimated(444) xor estimated(445);
partial_sums(2)(124) <= estimated(124) xor estimated(125);
partial_sums(2)(125) <= estimated(380) xor estimated(381);
partial_sums(2)(126) <= estimated(252) xor estimated(253);
partial_sums(2)(127) <= estimated(508) xor estimated(509);
partial_sums(2)(128) <= estimated(1);
partial_sums(2)(129) <= estimated(257);
partial_sums(2)(130) <= estimated(129);
partial_sums(2)(131) <= estimated(385);
partial_sums(2)(132) <= estimated(65);
partial_sums(2)(133) <= estimated(321);
partial_sums(2)(134) <= estimated(193);
partial_sums(2)(135) <= estimated(449);
partial_sums(2)(136) <= estimated(33);
partial_sums(2)(137) <= estimated(289);
partial_sums(2)(138) <= estimated(161);
partial_sums(2)(139) <= estimated(417);
partial_sums(2)(140) <= estimated(97);
partial_sums(2)(141) <= estimated(353);
partial_sums(2)(142) <= estimated(225);
partial_sums(2)(143) <= estimated(481);
partial_sums(2)(144) <= estimated(17);
partial_sums(2)(145) <= estimated(273);
partial_sums(2)(146) <= estimated(145);
partial_sums(2)(147) <= estimated(401);
partial_sums(2)(148) <= estimated(81);
partial_sums(2)(149) <= estimated(337);
partial_sums(2)(150) <= estimated(209);
partial_sums(2)(151) <= estimated(465);
partial_sums(2)(152) <= estimated(49);
partial_sums(2)(153) <= estimated(305);
partial_sums(2)(154) <= estimated(177);
partial_sums(2)(155) <= estimated(433);
partial_sums(2)(156) <= estimated(113);
partial_sums(2)(157) <= estimated(369);
partial_sums(2)(158) <= estimated(241);
partial_sums(2)(159) <= estimated(497);
partial_sums(2)(160) <= estimated(9);
partial_sums(2)(161) <= estimated(265);
partial_sums(2)(162) <= estimated(137);
partial_sums(2)(163) <= estimated(393);
partial_sums(2)(164) <= estimated(73);
partial_sums(2)(165) <= estimated(329);
partial_sums(2)(166) <= estimated(201);
partial_sums(2)(167) <= estimated(457);
partial_sums(2)(168) <= estimated(41);
partial_sums(2)(169) <= estimated(297);
partial_sums(2)(170) <= estimated(169);
partial_sums(2)(171) <= estimated(425);
partial_sums(2)(172) <= estimated(105);
partial_sums(2)(173) <= estimated(361);
partial_sums(2)(174) <= estimated(233);
partial_sums(2)(175) <= estimated(489);
partial_sums(2)(176) <= estimated(25);
partial_sums(2)(177) <= estimated(281);
partial_sums(2)(178) <= estimated(153);
partial_sums(2)(179) <= estimated(409);
partial_sums(2)(180) <= estimated(89);
partial_sums(2)(181) <= estimated(345);
partial_sums(2)(182) <= estimated(217);
partial_sums(2)(183) <= estimated(473);
partial_sums(2)(184) <= estimated(57);
partial_sums(2)(185) <= estimated(313);
partial_sums(2)(186) <= estimated(185);
partial_sums(2)(187) <= estimated(441);
partial_sums(2)(188) <= estimated(121);
partial_sums(2)(189) <= estimated(377);
partial_sums(2)(190) <= estimated(249);
partial_sums(2)(191) <= estimated(505);
partial_sums(2)(192) <= estimated(5);
partial_sums(2)(193) <= estimated(261);
partial_sums(2)(194) <= estimated(133);
partial_sums(2)(195) <= estimated(389);
partial_sums(2)(196) <= estimated(69);
partial_sums(2)(197) <= estimated(325);
partial_sums(2)(198) <= estimated(197);
partial_sums(2)(199) <= estimated(453);
partial_sums(2)(200) <= estimated(37);
partial_sums(2)(201) <= estimated(293);
partial_sums(2)(202) <= estimated(165);
partial_sums(2)(203) <= estimated(421);
partial_sums(2)(204) <= estimated(101);
partial_sums(2)(205) <= estimated(357);
partial_sums(2)(206) <= estimated(229);
partial_sums(2)(207) <= estimated(485);
partial_sums(2)(208) <= estimated(21);
partial_sums(2)(209) <= estimated(277);
partial_sums(2)(210) <= estimated(149);
partial_sums(2)(211) <= estimated(405);
partial_sums(2)(212) <= estimated(85);
partial_sums(2)(213) <= estimated(341);
partial_sums(2)(214) <= estimated(213);
partial_sums(2)(215) <= estimated(469);
partial_sums(2)(216) <= estimated(53);
partial_sums(2)(217) <= estimated(309);
partial_sums(2)(218) <= estimated(181);
partial_sums(2)(219) <= estimated(437);
partial_sums(2)(220) <= estimated(117);
partial_sums(2)(221) <= estimated(373);
partial_sums(2)(222) <= estimated(245);
partial_sums(2)(223) <= estimated(501);
partial_sums(2)(224) <= estimated(13);
partial_sums(2)(225) <= estimated(269);
partial_sums(2)(226) <= estimated(141);
partial_sums(2)(227) <= estimated(397);
partial_sums(2)(228) <= estimated(77);
partial_sums(2)(229) <= estimated(333);
partial_sums(2)(230) <= estimated(205);
partial_sums(2)(231) <= estimated(461);
partial_sums(2)(232) <= estimated(45);
partial_sums(2)(233) <= estimated(301);
partial_sums(2)(234) <= estimated(173);
partial_sums(2)(235) <= estimated(429);
partial_sums(2)(236) <= estimated(109);
partial_sums(2)(237) <= estimated(365);
partial_sums(2)(238) <= estimated(237);
partial_sums(2)(239) <= estimated(493);
partial_sums(2)(240) <= estimated(29);
partial_sums(2)(241) <= estimated(285);
partial_sums(2)(242) <= estimated(157);
partial_sums(2)(243) <= estimated(413);
partial_sums(2)(244) <= estimated(93);
partial_sums(2)(245) <= estimated(349);
partial_sums(2)(246) <= estimated(221);
partial_sums(2)(247) <= estimated(477);
partial_sums(2)(248) <= estimated(61);
partial_sums(2)(249) <= estimated(317);
partial_sums(2)(250) <= estimated(189);
partial_sums(2)(251) <= estimated(445);
partial_sums(2)(252) <= estimated(125);
partial_sums(2)(253) <= estimated(381);
partial_sums(2)(254) <= estimated(253);
partial_sums(2)(255) <= estimated(509);
partial_sums(3)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3);
partial_sums(3)(1) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259);
partial_sums(3)(2) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131);
partial_sums(3)(3) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387);
partial_sums(3)(4) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67);
partial_sums(3)(5) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323);
partial_sums(3)(6) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195);
partial_sums(3)(7) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451);
partial_sums(3)(8) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35);
partial_sums(3)(9) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291);
partial_sums(3)(10) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163);
partial_sums(3)(11) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419);
partial_sums(3)(12) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99);
partial_sums(3)(13) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355);
partial_sums(3)(14) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227);
partial_sums(3)(15) <= estimated(480) xor estimated(481) xor estimated(482) xor estimated(483);
partial_sums(3)(16) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19);
partial_sums(3)(17) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275);
partial_sums(3)(18) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147);
partial_sums(3)(19) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403);
partial_sums(3)(20) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83);
partial_sums(3)(21) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339);
partial_sums(3)(22) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211);
partial_sums(3)(23) <= estimated(464) xor estimated(465) xor estimated(466) xor estimated(467);
partial_sums(3)(24) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51);
partial_sums(3)(25) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307);
partial_sums(3)(26) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179);
partial_sums(3)(27) <= estimated(432) xor estimated(433) xor estimated(434) xor estimated(435);
partial_sums(3)(28) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115);
partial_sums(3)(29) <= estimated(368) xor estimated(369) xor estimated(370) xor estimated(371);
partial_sums(3)(30) <= estimated(240) xor estimated(241) xor estimated(242) xor estimated(243);
partial_sums(3)(31) <= estimated(496) xor estimated(497) xor estimated(498) xor estimated(499);
partial_sums(3)(32) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11);
partial_sums(3)(33) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267);
partial_sums(3)(34) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139);
partial_sums(3)(35) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395);
partial_sums(3)(36) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75);
partial_sums(3)(37) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331);
partial_sums(3)(38) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203);
partial_sums(3)(39) <= estimated(456) xor estimated(457) xor estimated(458) xor estimated(459);
partial_sums(3)(40) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43);
partial_sums(3)(41) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299);
partial_sums(3)(42) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171);
partial_sums(3)(43) <= estimated(424) xor estimated(425) xor estimated(426) xor estimated(427);
partial_sums(3)(44) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107);
partial_sums(3)(45) <= estimated(360) xor estimated(361) xor estimated(362) xor estimated(363);
partial_sums(3)(46) <= estimated(232) xor estimated(233) xor estimated(234) xor estimated(235);
partial_sums(3)(47) <= estimated(488) xor estimated(489) xor estimated(490) xor estimated(491);
partial_sums(3)(48) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27);
partial_sums(3)(49) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283);
partial_sums(3)(50) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155);
partial_sums(3)(51) <= estimated(408) xor estimated(409) xor estimated(410) xor estimated(411);
partial_sums(3)(52) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91);
partial_sums(3)(53) <= estimated(344) xor estimated(345) xor estimated(346) xor estimated(347);
partial_sums(3)(54) <= estimated(216) xor estimated(217) xor estimated(218) xor estimated(219);
partial_sums(3)(55) <= estimated(472) xor estimated(473) xor estimated(474) xor estimated(475);
partial_sums(3)(56) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59);
partial_sums(3)(57) <= estimated(312) xor estimated(313) xor estimated(314) xor estimated(315);
partial_sums(3)(58) <= estimated(184) xor estimated(185) xor estimated(186) xor estimated(187);
partial_sums(3)(59) <= estimated(440) xor estimated(441) xor estimated(442) xor estimated(443);
partial_sums(3)(60) <= estimated(120) xor estimated(121) xor estimated(122) xor estimated(123);
partial_sums(3)(61) <= estimated(376) xor estimated(377) xor estimated(378) xor estimated(379);
partial_sums(3)(62) <= estimated(248) xor estimated(249) xor estimated(250) xor estimated(251);
partial_sums(3)(63) <= estimated(504) xor estimated(505) xor estimated(506) xor estimated(507);
partial_sums(3)(64) <= estimated(2) xor estimated(3);
partial_sums(3)(65) <= estimated(258) xor estimated(259);
partial_sums(3)(66) <= estimated(130) xor estimated(131);
partial_sums(3)(67) <= estimated(386) xor estimated(387);
partial_sums(3)(68) <= estimated(66) xor estimated(67);
partial_sums(3)(69) <= estimated(322) xor estimated(323);
partial_sums(3)(70) <= estimated(194) xor estimated(195);
partial_sums(3)(71) <= estimated(450) xor estimated(451);
partial_sums(3)(72) <= estimated(34) xor estimated(35);
partial_sums(3)(73) <= estimated(290) xor estimated(291);
partial_sums(3)(74) <= estimated(162) xor estimated(163);
partial_sums(3)(75) <= estimated(418) xor estimated(419);
partial_sums(3)(76) <= estimated(98) xor estimated(99);
partial_sums(3)(77) <= estimated(354) xor estimated(355);
partial_sums(3)(78) <= estimated(226) xor estimated(227);
partial_sums(3)(79) <= estimated(482) xor estimated(483);
partial_sums(3)(80) <= estimated(18) xor estimated(19);
partial_sums(3)(81) <= estimated(274) xor estimated(275);
partial_sums(3)(82) <= estimated(146) xor estimated(147);
partial_sums(3)(83) <= estimated(402) xor estimated(403);
partial_sums(3)(84) <= estimated(82) xor estimated(83);
partial_sums(3)(85) <= estimated(338) xor estimated(339);
partial_sums(3)(86) <= estimated(210) xor estimated(211);
partial_sums(3)(87) <= estimated(466) xor estimated(467);
partial_sums(3)(88) <= estimated(50) xor estimated(51);
partial_sums(3)(89) <= estimated(306) xor estimated(307);
partial_sums(3)(90) <= estimated(178) xor estimated(179);
partial_sums(3)(91) <= estimated(434) xor estimated(435);
partial_sums(3)(92) <= estimated(114) xor estimated(115);
partial_sums(3)(93) <= estimated(370) xor estimated(371);
partial_sums(3)(94) <= estimated(242) xor estimated(243);
partial_sums(3)(95) <= estimated(498) xor estimated(499);
partial_sums(3)(96) <= estimated(10) xor estimated(11);
partial_sums(3)(97) <= estimated(266) xor estimated(267);
partial_sums(3)(98) <= estimated(138) xor estimated(139);
partial_sums(3)(99) <= estimated(394) xor estimated(395);
partial_sums(3)(100) <= estimated(74) xor estimated(75);
partial_sums(3)(101) <= estimated(330) xor estimated(331);
partial_sums(3)(102) <= estimated(202) xor estimated(203);
partial_sums(3)(103) <= estimated(458) xor estimated(459);
partial_sums(3)(104) <= estimated(42) xor estimated(43);
partial_sums(3)(105) <= estimated(298) xor estimated(299);
partial_sums(3)(106) <= estimated(170) xor estimated(171);
partial_sums(3)(107) <= estimated(426) xor estimated(427);
partial_sums(3)(108) <= estimated(106) xor estimated(107);
partial_sums(3)(109) <= estimated(362) xor estimated(363);
partial_sums(3)(110) <= estimated(234) xor estimated(235);
partial_sums(3)(111) <= estimated(490) xor estimated(491);
partial_sums(3)(112) <= estimated(26) xor estimated(27);
partial_sums(3)(113) <= estimated(282) xor estimated(283);
partial_sums(3)(114) <= estimated(154) xor estimated(155);
partial_sums(3)(115) <= estimated(410) xor estimated(411);
partial_sums(3)(116) <= estimated(90) xor estimated(91);
partial_sums(3)(117) <= estimated(346) xor estimated(347);
partial_sums(3)(118) <= estimated(218) xor estimated(219);
partial_sums(3)(119) <= estimated(474) xor estimated(475);
partial_sums(3)(120) <= estimated(58) xor estimated(59);
partial_sums(3)(121) <= estimated(314) xor estimated(315);
partial_sums(3)(122) <= estimated(186) xor estimated(187);
partial_sums(3)(123) <= estimated(442) xor estimated(443);
partial_sums(3)(124) <= estimated(122) xor estimated(123);
partial_sums(3)(125) <= estimated(378) xor estimated(379);
partial_sums(3)(126) <= estimated(250) xor estimated(251);
partial_sums(3)(127) <= estimated(506) xor estimated(507);
partial_sums(3)(128) <= estimated(1) xor estimated(3);
partial_sums(3)(129) <= estimated(257) xor estimated(259);
partial_sums(3)(130) <= estimated(129) xor estimated(131);
partial_sums(3)(131) <= estimated(385) xor estimated(387);
partial_sums(3)(132) <= estimated(65) xor estimated(67);
partial_sums(3)(133) <= estimated(321) xor estimated(323);
partial_sums(3)(134) <= estimated(193) xor estimated(195);
partial_sums(3)(135) <= estimated(449) xor estimated(451);
partial_sums(3)(136) <= estimated(33) xor estimated(35);
partial_sums(3)(137) <= estimated(289) xor estimated(291);
partial_sums(3)(138) <= estimated(161) xor estimated(163);
partial_sums(3)(139) <= estimated(417) xor estimated(419);
partial_sums(3)(140) <= estimated(97) xor estimated(99);
partial_sums(3)(141) <= estimated(353) xor estimated(355);
partial_sums(3)(142) <= estimated(225) xor estimated(227);
partial_sums(3)(143) <= estimated(481) xor estimated(483);
partial_sums(3)(144) <= estimated(17) xor estimated(19);
partial_sums(3)(145) <= estimated(273) xor estimated(275);
partial_sums(3)(146) <= estimated(145) xor estimated(147);
partial_sums(3)(147) <= estimated(401) xor estimated(403);
partial_sums(3)(148) <= estimated(81) xor estimated(83);
partial_sums(3)(149) <= estimated(337) xor estimated(339);
partial_sums(3)(150) <= estimated(209) xor estimated(211);
partial_sums(3)(151) <= estimated(465) xor estimated(467);
partial_sums(3)(152) <= estimated(49) xor estimated(51);
partial_sums(3)(153) <= estimated(305) xor estimated(307);
partial_sums(3)(154) <= estimated(177) xor estimated(179);
partial_sums(3)(155) <= estimated(433) xor estimated(435);
partial_sums(3)(156) <= estimated(113) xor estimated(115);
partial_sums(3)(157) <= estimated(369) xor estimated(371);
partial_sums(3)(158) <= estimated(241) xor estimated(243);
partial_sums(3)(159) <= estimated(497) xor estimated(499);
partial_sums(3)(160) <= estimated(9) xor estimated(11);
partial_sums(3)(161) <= estimated(265) xor estimated(267);
partial_sums(3)(162) <= estimated(137) xor estimated(139);
partial_sums(3)(163) <= estimated(393) xor estimated(395);
partial_sums(3)(164) <= estimated(73) xor estimated(75);
partial_sums(3)(165) <= estimated(329) xor estimated(331);
partial_sums(3)(166) <= estimated(201) xor estimated(203);
partial_sums(3)(167) <= estimated(457) xor estimated(459);
partial_sums(3)(168) <= estimated(41) xor estimated(43);
partial_sums(3)(169) <= estimated(297) xor estimated(299);
partial_sums(3)(170) <= estimated(169) xor estimated(171);
partial_sums(3)(171) <= estimated(425) xor estimated(427);
partial_sums(3)(172) <= estimated(105) xor estimated(107);
partial_sums(3)(173) <= estimated(361) xor estimated(363);
partial_sums(3)(174) <= estimated(233) xor estimated(235);
partial_sums(3)(175) <= estimated(489) xor estimated(491);
partial_sums(3)(176) <= estimated(25) xor estimated(27);
partial_sums(3)(177) <= estimated(281) xor estimated(283);
partial_sums(3)(178) <= estimated(153) xor estimated(155);
partial_sums(3)(179) <= estimated(409) xor estimated(411);
partial_sums(3)(180) <= estimated(89) xor estimated(91);
partial_sums(3)(181) <= estimated(345) xor estimated(347);
partial_sums(3)(182) <= estimated(217) xor estimated(219);
partial_sums(3)(183) <= estimated(473) xor estimated(475);
partial_sums(3)(184) <= estimated(57) xor estimated(59);
partial_sums(3)(185) <= estimated(313) xor estimated(315);
partial_sums(3)(186) <= estimated(185) xor estimated(187);
partial_sums(3)(187) <= estimated(441) xor estimated(443);
partial_sums(3)(188) <= estimated(121) xor estimated(123);
partial_sums(3)(189) <= estimated(377) xor estimated(379);
partial_sums(3)(190) <= estimated(249) xor estimated(251);
partial_sums(3)(191) <= estimated(505) xor estimated(507);
partial_sums(3)(192) <= estimated(3);
partial_sums(3)(193) <= estimated(259);
partial_sums(3)(194) <= estimated(131);
partial_sums(3)(195) <= estimated(387);
partial_sums(3)(196) <= estimated(67);
partial_sums(3)(197) <= estimated(323);
partial_sums(3)(198) <= estimated(195);
partial_sums(3)(199) <= estimated(451);
partial_sums(3)(200) <= estimated(35);
partial_sums(3)(201) <= estimated(291);
partial_sums(3)(202) <= estimated(163);
partial_sums(3)(203) <= estimated(419);
partial_sums(3)(204) <= estimated(99);
partial_sums(3)(205) <= estimated(355);
partial_sums(3)(206) <= estimated(227);
partial_sums(3)(207) <= estimated(483);
partial_sums(3)(208) <= estimated(19);
partial_sums(3)(209) <= estimated(275);
partial_sums(3)(210) <= estimated(147);
partial_sums(3)(211) <= estimated(403);
partial_sums(3)(212) <= estimated(83);
partial_sums(3)(213) <= estimated(339);
partial_sums(3)(214) <= estimated(211);
partial_sums(3)(215) <= estimated(467);
partial_sums(3)(216) <= estimated(51);
partial_sums(3)(217) <= estimated(307);
partial_sums(3)(218) <= estimated(179);
partial_sums(3)(219) <= estimated(435);
partial_sums(3)(220) <= estimated(115);
partial_sums(3)(221) <= estimated(371);
partial_sums(3)(222) <= estimated(243);
partial_sums(3)(223) <= estimated(499);
partial_sums(3)(224) <= estimated(11);
partial_sums(3)(225) <= estimated(267);
partial_sums(3)(226) <= estimated(139);
partial_sums(3)(227) <= estimated(395);
partial_sums(3)(228) <= estimated(75);
partial_sums(3)(229) <= estimated(331);
partial_sums(3)(230) <= estimated(203);
partial_sums(3)(231) <= estimated(459);
partial_sums(3)(232) <= estimated(43);
partial_sums(3)(233) <= estimated(299);
partial_sums(3)(234) <= estimated(171);
partial_sums(3)(235) <= estimated(427);
partial_sums(3)(236) <= estimated(107);
partial_sums(3)(237) <= estimated(363);
partial_sums(3)(238) <= estimated(235);
partial_sums(3)(239) <= estimated(491);
partial_sums(3)(240) <= estimated(27);
partial_sums(3)(241) <= estimated(283);
partial_sums(3)(242) <= estimated(155);
partial_sums(3)(243) <= estimated(411);
partial_sums(3)(244) <= estimated(91);
partial_sums(3)(245) <= estimated(347);
partial_sums(3)(246) <= estimated(219);
partial_sums(3)(247) <= estimated(475);
partial_sums(3)(248) <= estimated(59);
partial_sums(3)(249) <= estimated(315);
partial_sums(3)(250) <= estimated(187);
partial_sums(3)(251) <= estimated(443);
partial_sums(3)(252) <= estimated(123);
partial_sums(3)(253) <= estimated(379);
partial_sums(3)(254) <= estimated(251);
partial_sums(3)(255) <= estimated(507);
partial_sums(4)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7);
partial_sums(4)(1) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263);
partial_sums(4)(2) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135);
partial_sums(4)(3) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391);
partial_sums(4)(4) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71);
partial_sums(4)(5) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327);
partial_sums(4)(6) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199);
partial_sums(4)(7) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455);
partial_sums(4)(8) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39);
partial_sums(4)(9) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295);
partial_sums(4)(10) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167);
partial_sums(4)(11) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423);
partial_sums(4)(12) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103);
partial_sums(4)(13) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359);
partial_sums(4)(14) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231);
partial_sums(4)(15) <= estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487);
partial_sums(4)(16) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23);
partial_sums(4)(17) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279);
partial_sums(4)(18) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151);
partial_sums(4)(19) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407);
partial_sums(4)(20) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87);
partial_sums(4)(21) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343);
partial_sums(4)(22) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215);
partial_sums(4)(23) <= estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471);
partial_sums(4)(24) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55);
partial_sums(4)(25) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311);
partial_sums(4)(26) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183);
partial_sums(4)(27) <= estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439);
partial_sums(4)(28) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119);
partial_sums(4)(29) <= estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375);
partial_sums(4)(30) <= estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247);
partial_sums(4)(31) <= estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503);
partial_sums(4)(32) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7);
partial_sums(4)(33) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263);
partial_sums(4)(34) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135);
partial_sums(4)(35) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391);
partial_sums(4)(36) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71);
partial_sums(4)(37) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327);
partial_sums(4)(38) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199);
partial_sums(4)(39) <= estimated(452) xor estimated(453) xor estimated(454) xor estimated(455);
partial_sums(4)(40) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39);
partial_sums(4)(41) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295);
partial_sums(4)(42) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167);
partial_sums(4)(43) <= estimated(420) xor estimated(421) xor estimated(422) xor estimated(423);
partial_sums(4)(44) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103);
partial_sums(4)(45) <= estimated(356) xor estimated(357) xor estimated(358) xor estimated(359);
partial_sums(4)(46) <= estimated(228) xor estimated(229) xor estimated(230) xor estimated(231);
partial_sums(4)(47) <= estimated(484) xor estimated(485) xor estimated(486) xor estimated(487);
partial_sums(4)(48) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23);
partial_sums(4)(49) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279);
partial_sums(4)(50) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151);
partial_sums(4)(51) <= estimated(404) xor estimated(405) xor estimated(406) xor estimated(407);
partial_sums(4)(52) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87);
partial_sums(4)(53) <= estimated(340) xor estimated(341) xor estimated(342) xor estimated(343);
partial_sums(4)(54) <= estimated(212) xor estimated(213) xor estimated(214) xor estimated(215);
partial_sums(4)(55) <= estimated(468) xor estimated(469) xor estimated(470) xor estimated(471);
partial_sums(4)(56) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55);
partial_sums(4)(57) <= estimated(308) xor estimated(309) xor estimated(310) xor estimated(311);
partial_sums(4)(58) <= estimated(180) xor estimated(181) xor estimated(182) xor estimated(183);
partial_sums(4)(59) <= estimated(436) xor estimated(437) xor estimated(438) xor estimated(439);
partial_sums(4)(60) <= estimated(116) xor estimated(117) xor estimated(118) xor estimated(119);
partial_sums(4)(61) <= estimated(372) xor estimated(373) xor estimated(374) xor estimated(375);
partial_sums(4)(62) <= estimated(244) xor estimated(245) xor estimated(246) xor estimated(247);
partial_sums(4)(63) <= estimated(500) xor estimated(501) xor estimated(502) xor estimated(503);
partial_sums(4)(64) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7);
partial_sums(4)(65) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263);
partial_sums(4)(66) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135);
partial_sums(4)(67) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391);
partial_sums(4)(68) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71);
partial_sums(4)(69) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327);
partial_sums(4)(70) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199);
partial_sums(4)(71) <= estimated(450) xor estimated(451) xor estimated(454) xor estimated(455);
partial_sums(4)(72) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39);
partial_sums(4)(73) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295);
partial_sums(4)(74) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167);
partial_sums(4)(75) <= estimated(418) xor estimated(419) xor estimated(422) xor estimated(423);
partial_sums(4)(76) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103);
partial_sums(4)(77) <= estimated(354) xor estimated(355) xor estimated(358) xor estimated(359);
partial_sums(4)(78) <= estimated(226) xor estimated(227) xor estimated(230) xor estimated(231);
partial_sums(4)(79) <= estimated(482) xor estimated(483) xor estimated(486) xor estimated(487);
partial_sums(4)(80) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23);
partial_sums(4)(81) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279);
partial_sums(4)(82) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151);
partial_sums(4)(83) <= estimated(402) xor estimated(403) xor estimated(406) xor estimated(407);
partial_sums(4)(84) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87);
partial_sums(4)(85) <= estimated(338) xor estimated(339) xor estimated(342) xor estimated(343);
partial_sums(4)(86) <= estimated(210) xor estimated(211) xor estimated(214) xor estimated(215);
partial_sums(4)(87) <= estimated(466) xor estimated(467) xor estimated(470) xor estimated(471);
partial_sums(4)(88) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55);
partial_sums(4)(89) <= estimated(306) xor estimated(307) xor estimated(310) xor estimated(311);
partial_sums(4)(90) <= estimated(178) xor estimated(179) xor estimated(182) xor estimated(183);
partial_sums(4)(91) <= estimated(434) xor estimated(435) xor estimated(438) xor estimated(439);
partial_sums(4)(92) <= estimated(114) xor estimated(115) xor estimated(118) xor estimated(119);
partial_sums(4)(93) <= estimated(370) xor estimated(371) xor estimated(374) xor estimated(375);
partial_sums(4)(94) <= estimated(242) xor estimated(243) xor estimated(246) xor estimated(247);
partial_sums(4)(95) <= estimated(498) xor estimated(499) xor estimated(502) xor estimated(503);
partial_sums(4)(96) <= estimated(6) xor estimated(7);
partial_sums(4)(97) <= estimated(262) xor estimated(263);
partial_sums(4)(98) <= estimated(134) xor estimated(135);
partial_sums(4)(99) <= estimated(390) xor estimated(391);
partial_sums(4)(100) <= estimated(70) xor estimated(71);
partial_sums(4)(101) <= estimated(326) xor estimated(327);
partial_sums(4)(102) <= estimated(198) xor estimated(199);
partial_sums(4)(103) <= estimated(454) xor estimated(455);
partial_sums(4)(104) <= estimated(38) xor estimated(39);
partial_sums(4)(105) <= estimated(294) xor estimated(295);
partial_sums(4)(106) <= estimated(166) xor estimated(167);
partial_sums(4)(107) <= estimated(422) xor estimated(423);
partial_sums(4)(108) <= estimated(102) xor estimated(103);
partial_sums(4)(109) <= estimated(358) xor estimated(359);
partial_sums(4)(110) <= estimated(230) xor estimated(231);
partial_sums(4)(111) <= estimated(486) xor estimated(487);
partial_sums(4)(112) <= estimated(22) xor estimated(23);
partial_sums(4)(113) <= estimated(278) xor estimated(279);
partial_sums(4)(114) <= estimated(150) xor estimated(151);
partial_sums(4)(115) <= estimated(406) xor estimated(407);
partial_sums(4)(116) <= estimated(86) xor estimated(87);
partial_sums(4)(117) <= estimated(342) xor estimated(343);
partial_sums(4)(118) <= estimated(214) xor estimated(215);
partial_sums(4)(119) <= estimated(470) xor estimated(471);
partial_sums(4)(120) <= estimated(54) xor estimated(55);
partial_sums(4)(121) <= estimated(310) xor estimated(311);
partial_sums(4)(122) <= estimated(182) xor estimated(183);
partial_sums(4)(123) <= estimated(438) xor estimated(439);
partial_sums(4)(124) <= estimated(118) xor estimated(119);
partial_sums(4)(125) <= estimated(374) xor estimated(375);
partial_sums(4)(126) <= estimated(246) xor estimated(247);
partial_sums(4)(127) <= estimated(502) xor estimated(503);
partial_sums(4)(128) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7);
partial_sums(4)(129) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263);
partial_sums(4)(130) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135);
partial_sums(4)(131) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391);
partial_sums(4)(132) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71);
partial_sums(4)(133) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327);
partial_sums(4)(134) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199);
partial_sums(4)(135) <= estimated(449) xor estimated(451) xor estimated(453) xor estimated(455);
partial_sums(4)(136) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39);
partial_sums(4)(137) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295);
partial_sums(4)(138) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167);
partial_sums(4)(139) <= estimated(417) xor estimated(419) xor estimated(421) xor estimated(423);
partial_sums(4)(140) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103);
partial_sums(4)(141) <= estimated(353) xor estimated(355) xor estimated(357) xor estimated(359);
partial_sums(4)(142) <= estimated(225) xor estimated(227) xor estimated(229) xor estimated(231);
partial_sums(4)(143) <= estimated(481) xor estimated(483) xor estimated(485) xor estimated(487);
partial_sums(4)(144) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23);
partial_sums(4)(145) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279);
partial_sums(4)(146) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151);
partial_sums(4)(147) <= estimated(401) xor estimated(403) xor estimated(405) xor estimated(407);
partial_sums(4)(148) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87);
partial_sums(4)(149) <= estimated(337) xor estimated(339) xor estimated(341) xor estimated(343);
partial_sums(4)(150) <= estimated(209) xor estimated(211) xor estimated(213) xor estimated(215);
partial_sums(4)(151) <= estimated(465) xor estimated(467) xor estimated(469) xor estimated(471);
partial_sums(4)(152) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55);
partial_sums(4)(153) <= estimated(305) xor estimated(307) xor estimated(309) xor estimated(311);
partial_sums(4)(154) <= estimated(177) xor estimated(179) xor estimated(181) xor estimated(183);
partial_sums(4)(155) <= estimated(433) xor estimated(435) xor estimated(437) xor estimated(439);
partial_sums(4)(156) <= estimated(113) xor estimated(115) xor estimated(117) xor estimated(119);
partial_sums(4)(157) <= estimated(369) xor estimated(371) xor estimated(373) xor estimated(375);
partial_sums(4)(158) <= estimated(241) xor estimated(243) xor estimated(245) xor estimated(247);
partial_sums(4)(159) <= estimated(497) xor estimated(499) xor estimated(501) xor estimated(503);
partial_sums(4)(160) <= estimated(5) xor estimated(7);
partial_sums(4)(161) <= estimated(261) xor estimated(263);
partial_sums(4)(162) <= estimated(133) xor estimated(135);
partial_sums(4)(163) <= estimated(389) xor estimated(391);
partial_sums(4)(164) <= estimated(69) xor estimated(71);
partial_sums(4)(165) <= estimated(325) xor estimated(327);
partial_sums(4)(166) <= estimated(197) xor estimated(199);
partial_sums(4)(167) <= estimated(453) xor estimated(455);
partial_sums(4)(168) <= estimated(37) xor estimated(39);
partial_sums(4)(169) <= estimated(293) xor estimated(295);
partial_sums(4)(170) <= estimated(165) xor estimated(167);
partial_sums(4)(171) <= estimated(421) xor estimated(423);
partial_sums(4)(172) <= estimated(101) xor estimated(103);
partial_sums(4)(173) <= estimated(357) xor estimated(359);
partial_sums(4)(174) <= estimated(229) xor estimated(231);
partial_sums(4)(175) <= estimated(485) xor estimated(487);
partial_sums(4)(176) <= estimated(21) xor estimated(23);
partial_sums(4)(177) <= estimated(277) xor estimated(279);
partial_sums(4)(178) <= estimated(149) xor estimated(151);
partial_sums(4)(179) <= estimated(405) xor estimated(407);
partial_sums(4)(180) <= estimated(85) xor estimated(87);
partial_sums(4)(181) <= estimated(341) xor estimated(343);
partial_sums(4)(182) <= estimated(213) xor estimated(215);
partial_sums(4)(183) <= estimated(469) xor estimated(471);
partial_sums(4)(184) <= estimated(53) xor estimated(55);
partial_sums(4)(185) <= estimated(309) xor estimated(311);
partial_sums(4)(186) <= estimated(181) xor estimated(183);
partial_sums(4)(187) <= estimated(437) xor estimated(439);
partial_sums(4)(188) <= estimated(117) xor estimated(119);
partial_sums(4)(189) <= estimated(373) xor estimated(375);
partial_sums(4)(190) <= estimated(245) xor estimated(247);
partial_sums(4)(191) <= estimated(501) xor estimated(503);
partial_sums(4)(192) <= estimated(3) xor estimated(7);
partial_sums(4)(193) <= estimated(259) xor estimated(263);
partial_sums(4)(194) <= estimated(131) xor estimated(135);
partial_sums(4)(195) <= estimated(387) xor estimated(391);
partial_sums(4)(196) <= estimated(67) xor estimated(71);
partial_sums(4)(197) <= estimated(323) xor estimated(327);
partial_sums(4)(198) <= estimated(195) xor estimated(199);
partial_sums(4)(199) <= estimated(451) xor estimated(455);
partial_sums(4)(200) <= estimated(35) xor estimated(39);
partial_sums(4)(201) <= estimated(291) xor estimated(295);
partial_sums(4)(202) <= estimated(163) xor estimated(167);
partial_sums(4)(203) <= estimated(419) xor estimated(423);
partial_sums(4)(204) <= estimated(99) xor estimated(103);
partial_sums(4)(205) <= estimated(355) xor estimated(359);
partial_sums(4)(206) <= estimated(227) xor estimated(231);
partial_sums(4)(207) <= estimated(483) xor estimated(487);
partial_sums(4)(208) <= estimated(19) xor estimated(23);
partial_sums(4)(209) <= estimated(275) xor estimated(279);
partial_sums(4)(210) <= estimated(147) xor estimated(151);
partial_sums(4)(211) <= estimated(403) xor estimated(407);
partial_sums(4)(212) <= estimated(83) xor estimated(87);
partial_sums(4)(213) <= estimated(339) xor estimated(343);
partial_sums(4)(214) <= estimated(211) xor estimated(215);
partial_sums(4)(215) <= estimated(467) xor estimated(471);
partial_sums(4)(216) <= estimated(51) xor estimated(55);
partial_sums(4)(217) <= estimated(307) xor estimated(311);
partial_sums(4)(218) <= estimated(179) xor estimated(183);
partial_sums(4)(219) <= estimated(435) xor estimated(439);
partial_sums(4)(220) <= estimated(115) xor estimated(119);
partial_sums(4)(221) <= estimated(371) xor estimated(375);
partial_sums(4)(222) <= estimated(243) xor estimated(247);
partial_sums(4)(223) <= estimated(499) xor estimated(503);
partial_sums(4)(224) <= estimated(7);
partial_sums(4)(225) <= estimated(263);
partial_sums(4)(226) <= estimated(135);
partial_sums(4)(227) <= estimated(391);
partial_sums(4)(228) <= estimated(71);
partial_sums(4)(229) <= estimated(327);
partial_sums(4)(230) <= estimated(199);
partial_sums(4)(231) <= estimated(455);
partial_sums(4)(232) <= estimated(39);
partial_sums(4)(233) <= estimated(295);
partial_sums(4)(234) <= estimated(167);
partial_sums(4)(235) <= estimated(423);
partial_sums(4)(236) <= estimated(103);
partial_sums(4)(237) <= estimated(359);
partial_sums(4)(238) <= estimated(231);
partial_sums(4)(239) <= estimated(487);
partial_sums(4)(240) <= estimated(23);
partial_sums(4)(241) <= estimated(279);
partial_sums(4)(242) <= estimated(151);
partial_sums(4)(243) <= estimated(407);
partial_sums(4)(244) <= estimated(87);
partial_sums(4)(245) <= estimated(343);
partial_sums(4)(246) <= estimated(215);
partial_sums(4)(247) <= estimated(471);
partial_sums(4)(248) <= estimated(55);
partial_sums(4)(249) <= estimated(311);
partial_sums(4)(250) <= estimated(183);
partial_sums(4)(251) <= estimated(439);
partial_sums(4)(252) <= estimated(119);
partial_sums(4)(253) <= estimated(375);
partial_sums(4)(254) <= estimated(247);
partial_sums(4)(255) <= estimated(503);
partial_sums(5)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(1) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(2) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(3) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(4) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(5) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(6) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(7) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(8) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(9) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(10) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(11) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(12) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(13) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(14) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(15) <= estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(16) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(17) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(18) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(19) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(20) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(21) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(22) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(23) <= estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(24) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(25) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(26) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(27) <= estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(28) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(29) <= estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(30) <= estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(31) <= estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(32) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(33) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(34) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(35) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(36) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(37) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(38) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(39) <= estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(40) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(41) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(42) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(43) <= estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(44) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(45) <= estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(46) <= estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(47) <= estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(48) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(49) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(50) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(51) <= estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(52) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(53) <= estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(54) <= estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(55) <= estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(56) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(57) <= estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(58) <= estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(59) <= estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(60) <= estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(61) <= estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(62) <= estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(63) <= estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(64) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15);
partial_sums(5)(65) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271);
partial_sums(5)(66) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143);
partial_sums(5)(67) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399);
partial_sums(5)(68) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79);
partial_sums(5)(69) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335);
partial_sums(5)(70) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207);
partial_sums(5)(71) <= estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463);
partial_sums(5)(72) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47);
partial_sums(5)(73) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303);
partial_sums(5)(74) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175);
partial_sums(5)(75) <= estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431);
partial_sums(5)(76) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111);
partial_sums(5)(77) <= estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367);
partial_sums(5)(78) <= estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239);
partial_sums(5)(79) <= estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495);
partial_sums(5)(80) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15);
partial_sums(5)(81) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271);
partial_sums(5)(82) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143);
partial_sums(5)(83) <= estimated(394) xor estimated(395) xor estimated(398) xor estimated(399);
partial_sums(5)(84) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79);
partial_sums(5)(85) <= estimated(330) xor estimated(331) xor estimated(334) xor estimated(335);
partial_sums(5)(86) <= estimated(202) xor estimated(203) xor estimated(206) xor estimated(207);
partial_sums(5)(87) <= estimated(458) xor estimated(459) xor estimated(462) xor estimated(463);
partial_sums(5)(88) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47);
partial_sums(5)(89) <= estimated(298) xor estimated(299) xor estimated(302) xor estimated(303);
partial_sums(5)(90) <= estimated(170) xor estimated(171) xor estimated(174) xor estimated(175);
partial_sums(5)(91) <= estimated(426) xor estimated(427) xor estimated(430) xor estimated(431);
partial_sums(5)(92) <= estimated(106) xor estimated(107) xor estimated(110) xor estimated(111);
partial_sums(5)(93) <= estimated(362) xor estimated(363) xor estimated(366) xor estimated(367);
partial_sums(5)(94) <= estimated(234) xor estimated(235) xor estimated(238) xor estimated(239);
partial_sums(5)(95) <= estimated(490) xor estimated(491) xor estimated(494) xor estimated(495);
partial_sums(5)(96) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15);
partial_sums(5)(97) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271);
partial_sums(5)(98) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143);
partial_sums(5)(99) <= estimated(390) xor estimated(391) xor estimated(398) xor estimated(399);
partial_sums(5)(100) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79);
partial_sums(5)(101) <= estimated(326) xor estimated(327) xor estimated(334) xor estimated(335);
partial_sums(5)(102) <= estimated(198) xor estimated(199) xor estimated(206) xor estimated(207);
partial_sums(5)(103) <= estimated(454) xor estimated(455) xor estimated(462) xor estimated(463);
partial_sums(5)(104) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47);
partial_sums(5)(105) <= estimated(294) xor estimated(295) xor estimated(302) xor estimated(303);
partial_sums(5)(106) <= estimated(166) xor estimated(167) xor estimated(174) xor estimated(175);
partial_sums(5)(107) <= estimated(422) xor estimated(423) xor estimated(430) xor estimated(431);
partial_sums(5)(108) <= estimated(102) xor estimated(103) xor estimated(110) xor estimated(111);
partial_sums(5)(109) <= estimated(358) xor estimated(359) xor estimated(366) xor estimated(367);
partial_sums(5)(110) <= estimated(230) xor estimated(231) xor estimated(238) xor estimated(239);
partial_sums(5)(111) <= estimated(486) xor estimated(487) xor estimated(494) xor estimated(495);
partial_sums(5)(112) <= estimated(14) xor estimated(15);
partial_sums(5)(113) <= estimated(270) xor estimated(271);
partial_sums(5)(114) <= estimated(142) xor estimated(143);
partial_sums(5)(115) <= estimated(398) xor estimated(399);
partial_sums(5)(116) <= estimated(78) xor estimated(79);
partial_sums(5)(117) <= estimated(334) xor estimated(335);
partial_sums(5)(118) <= estimated(206) xor estimated(207);
partial_sums(5)(119) <= estimated(462) xor estimated(463);
partial_sums(5)(120) <= estimated(46) xor estimated(47);
partial_sums(5)(121) <= estimated(302) xor estimated(303);
partial_sums(5)(122) <= estimated(174) xor estimated(175);
partial_sums(5)(123) <= estimated(430) xor estimated(431);
partial_sums(5)(124) <= estimated(110) xor estimated(111);
partial_sums(5)(125) <= estimated(366) xor estimated(367);
partial_sums(5)(126) <= estimated(238) xor estimated(239);
partial_sums(5)(127) <= estimated(494) xor estimated(495);
partial_sums(5)(128) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15);
partial_sums(5)(129) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271);
partial_sums(5)(130) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143);
partial_sums(5)(131) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399);
partial_sums(5)(132) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79);
partial_sums(5)(133) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335);
partial_sums(5)(134) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207);
partial_sums(5)(135) <= estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463);
partial_sums(5)(136) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47);
partial_sums(5)(137) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303);
partial_sums(5)(138) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175);
partial_sums(5)(139) <= estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431);
partial_sums(5)(140) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111);
partial_sums(5)(141) <= estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367);
partial_sums(5)(142) <= estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239);
partial_sums(5)(143) <= estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495);
partial_sums(5)(144) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15);
partial_sums(5)(145) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271);
partial_sums(5)(146) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143);
partial_sums(5)(147) <= estimated(393) xor estimated(395) xor estimated(397) xor estimated(399);
partial_sums(5)(148) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79);
partial_sums(5)(149) <= estimated(329) xor estimated(331) xor estimated(333) xor estimated(335);
partial_sums(5)(150) <= estimated(201) xor estimated(203) xor estimated(205) xor estimated(207);
partial_sums(5)(151) <= estimated(457) xor estimated(459) xor estimated(461) xor estimated(463);
partial_sums(5)(152) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47);
partial_sums(5)(153) <= estimated(297) xor estimated(299) xor estimated(301) xor estimated(303);
partial_sums(5)(154) <= estimated(169) xor estimated(171) xor estimated(173) xor estimated(175);
partial_sums(5)(155) <= estimated(425) xor estimated(427) xor estimated(429) xor estimated(431);
partial_sums(5)(156) <= estimated(105) xor estimated(107) xor estimated(109) xor estimated(111);
partial_sums(5)(157) <= estimated(361) xor estimated(363) xor estimated(365) xor estimated(367);
partial_sums(5)(158) <= estimated(233) xor estimated(235) xor estimated(237) xor estimated(239);
partial_sums(5)(159) <= estimated(489) xor estimated(491) xor estimated(493) xor estimated(495);
partial_sums(5)(160) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15);
partial_sums(5)(161) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271);
partial_sums(5)(162) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143);
partial_sums(5)(163) <= estimated(389) xor estimated(391) xor estimated(397) xor estimated(399);
partial_sums(5)(164) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79);
partial_sums(5)(165) <= estimated(325) xor estimated(327) xor estimated(333) xor estimated(335);
partial_sums(5)(166) <= estimated(197) xor estimated(199) xor estimated(205) xor estimated(207);
partial_sums(5)(167) <= estimated(453) xor estimated(455) xor estimated(461) xor estimated(463);
partial_sums(5)(168) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47);
partial_sums(5)(169) <= estimated(293) xor estimated(295) xor estimated(301) xor estimated(303);
partial_sums(5)(170) <= estimated(165) xor estimated(167) xor estimated(173) xor estimated(175);
partial_sums(5)(171) <= estimated(421) xor estimated(423) xor estimated(429) xor estimated(431);
partial_sums(5)(172) <= estimated(101) xor estimated(103) xor estimated(109) xor estimated(111);
partial_sums(5)(173) <= estimated(357) xor estimated(359) xor estimated(365) xor estimated(367);
partial_sums(5)(174) <= estimated(229) xor estimated(231) xor estimated(237) xor estimated(239);
partial_sums(5)(175) <= estimated(485) xor estimated(487) xor estimated(493) xor estimated(495);
partial_sums(5)(176) <= estimated(13) xor estimated(15);
partial_sums(5)(177) <= estimated(269) xor estimated(271);
partial_sums(5)(178) <= estimated(141) xor estimated(143);
partial_sums(5)(179) <= estimated(397) xor estimated(399);
partial_sums(5)(180) <= estimated(77) xor estimated(79);
partial_sums(5)(181) <= estimated(333) xor estimated(335);
partial_sums(5)(182) <= estimated(205) xor estimated(207);
partial_sums(5)(183) <= estimated(461) xor estimated(463);
partial_sums(5)(184) <= estimated(45) xor estimated(47);
partial_sums(5)(185) <= estimated(301) xor estimated(303);
partial_sums(5)(186) <= estimated(173) xor estimated(175);
partial_sums(5)(187) <= estimated(429) xor estimated(431);
partial_sums(5)(188) <= estimated(109) xor estimated(111);
partial_sums(5)(189) <= estimated(365) xor estimated(367);
partial_sums(5)(190) <= estimated(237) xor estimated(239);
partial_sums(5)(191) <= estimated(493) xor estimated(495);
partial_sums(5)(192) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15);
partial_sums(5)(193) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271);
partial_sums(5)(194) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143);
partial_sums(5)(195) <= estimated(387) xor estimated(391) xor estimated(395) xor estimated(399);
partial_sums(5)(196) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79);
partial_sums(5)(197) <= estimated(323) xor estimated(327) xor estimated(331) xor estimated(335);
partial_sums(5)(198) <= estimated(195) xor estimated(199) xor estimated(203) xor estimated(207);
partial_sums(5)(199) <= estimated(451) xor estimated(455) xor estimated(459) xor estimated(463);
partial_sums(5)(200) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47);
partial_sums(5)(201) <= estimated(291) xor estimated(295) xor estimated(299) xor estimated(303);
partial_sums(5)(202) <= estimated(163) xor estimated(167) xor estimated(171) xor estimated(175);
partial_sums(5)(203) <= estimated(419) xor estimated(423) xor estimated(427) xor estimated(431);
partial_sums(5)(204) <= estimated(99) xor estimated(103) xor estimated(107) xor estimated(111);
partial_sums(5)(205) <= estimated(355) xor estimated(359) xor estimated(363) xor estimated(367);
partial_sums(5)(206) <= estimated(227) xor estimated(231) xor estimated(235) xor estimated(239);
partial_sums(5)(207) <= estimated(483) xor estimated(487) xor estimated(491) xor estimated(495);
partial_sums(5)(208) <= estimated(11) xor estimated(15);
partial_sums(5)(209) <= estimated(267) xor estimated(271);
partial_sums(5)(210) <= estimated(139) xor estimated(143);
partial_sums(5)(211) <= estimated(395) xor estimated(399);
partial_sums(5)(212) <= estimated(75) xor estimated(79);
partial_sums(5)(213) <= estimated(331) xor estimated(335);
partial_sums(5)(214) <= estimated(203) xor estimated(207);
partial_sums(5)(215) <= estimated(459) xor estimated(463);
partial_sums(5)(216) <= estimated(43) xor estimated(47);
partial_sums(5)(217) <= estimated(299) xor estimated(303);
partial_sums(5)(218) <= estimated(171) xor estimated(175);
partial_sums(5)(219) <= estimated(427) xor estimated(431);
partial_sums(5)(220) <= estimated(107) xor estimated(111);
partial_sums(5)(221) <= estimated(363) xor estimated(367);
partial_sums(5)(222) <= estimated(235) xor estimated(239);
partial_sums(5)(223) <= estimated(491) xor estimated(495);
partial_sums(5)(224) <= estimated(7) xor estimated(15);
partial_sums(5)(225) <= estimated(263) xor estimated(271);
partial_sums(5)(226) <= estimated(135) xor estimated(143);
partial_sums(5)(227) <= estimated(391) xor estimated(399);
partial_sums(5)(228) <= estimated(71) xor estimated(79);
partial_sums(5)(229) <= estimated(327) xor estimated(335);
partial_sums(5)(230) <= estimated(199) xor estimated(207);
partial_sums(5)(231) <= estimated(455) xor estimated(463);
partial_sums(5)(232) <= estimated(39) xor estimated(47);
partial_sums(5)(233) <= estimated(295) xor estimated(303);
partial_sums(5)(234) <= estimated(167) xor estimated(175);
partial_sums(5)(235) <= estimated(423) xor estimated(431);
partial_sums(5)(236) <= estimated(103) xor estimated(111);
partial_sums(5)(237) <= estimated(359) xor estimated(367);
partial_sums(5)(238) <= estimated(231) xor estimated(239);
partial_sums(5)(239) <= estimated(487) xor estimated(495);
partial_sums(5)(240) <= estimated(15);
partial_sums(5)(241) <= estimated(271);
partial_sums(5)(242) <= estimated(143);
partial_sums(5)(243) <= estimated(399);
partial_sums(5)(244) <= estimated(79);
partial_sums(5)(245) <= estimated(335);
partial_sums(5)(246) <= estimated(207);
partial_sums(5)(247) <= estimated(463);
partial_sums(5)(248) <= estimated(47);
partial_sums(5)(249) <= estimated(303);
partial_sums(5)(250) <= estimated(175);
partial_sums(5)(251) <= estimated(431);
partial_sums(5)(252) <= estimated(111);
partial_sums(5)(253) <= estimated(367);
partial_sums(5)(254) <= estimated(239);
partial_sums(5)(255) <= estimated(495);
partial_sums(6)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(1) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(2) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(3) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(4) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(5) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(6) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(7) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(8) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(9) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(10) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(11) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(12) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(13) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(14) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(15) <= estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(16) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(17) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(18) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(19) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(20) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(21) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(22) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(23) <= estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(24) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(25) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(26) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(27) <= estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(28) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(29) <= estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(30) <= estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(31) <= estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(32) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(33) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(34) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(35) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(36) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(37) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(38) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(39) <= estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(40) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(41) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(42) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(43) <= estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(44) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(45) <= estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(46) <= estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(47) <= estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(48) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(49) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(50) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(51) <= estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(52) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(53) <= estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(54) <= estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(55) <= estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(56) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(57) <= estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(58) <= estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(59) <= estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(60) <= estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(61) <= estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(62) <= estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(63) <= estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(64) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(65) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(66) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(67) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(68) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(69) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(70) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(71) <= estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(72) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(73) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(74) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(75) <= estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(76) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(77) <= estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(78) <= estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(79) <= estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(80) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(81) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(82) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(83) <= estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(84) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(85) <= estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(86) <= estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(87) <= estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(88) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(89) <= estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(90) <= estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(91) <= estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(92) <= estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(93) <= estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(94) <= estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(95) <= estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(96) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31);
partial_sums(6)(97) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287);
partial_sums(6)(98) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159);
partial_sums(6)(99) <= estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415);
partial_sums(6)(100) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95);
partial_sums(6)(101) <= estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351);
partial_sums(6)(102) <= estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223);
partial_sums(6)(103) <= estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479);
partial_sums(6)(104) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31);
partial_sums(6)(105) <= estimated(278) xor estimated(279) xor estimated(286) xor estimated(287);
partial_sums(6)(106) <= estimated(150) xor estimated(151) xor estimated(158) xor estimated(159);
partial_sums(6)(107) <= estimated(406) xor estimated(407) xor estimated(414) xor estimated(415);
partial_sums(6)(108) <= estimated(86) xor estimated(87) xor estimated(94) xor estimated(95);
partial_sums(6)(109) <= estimated(342) xor estimated(343) xor estimated(350) xor estimated(351);
partial_sums(6)(110) <= estimated(214) xor estimated(215) xor estimated(222) xor estimated(223);
partial_sums(6)(111) <= estimated(470) xor estimated(471) xor estimated(478) xor estimated(479);
partial_sums(6)(112) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31);
partial_sums(6)(113) <= estimated(270) xor estimated(271) xor estimated(286) xor estimated(287);
partial_sums(6)(114) <= estimated(142) xor estimated(143) xor estimated(158) xor estimated(159);
partial_sums(6)(115) <= estimated(398) xor estimated(399) xor estimated(414) xor estimated(415);
partial_sums(6)(116) <= estimated(78) xor estimated(79) xor estimated(94) xor estimated(95);
partial_sums(6)(117) <= estimated(334) xor estimated(335) xor estimated(350) xor estimated(351);
partial_sums(6)(118) <= estimated(206) xor estimated(207) xor estimated(222) xor estimated(223);
partial_sums(6)(119) <= estimated(462) xor estimated(463) xor estimated(478) xor estimated(479);
partial_sums(6)(120) <= estimated(30) xor estimated(31);
partial_sums(6)(121) <= estimated(286) xor estimated(287);
partial_sums(6)(122) <= estimated(158) xor estimated(159);
partial_sums(6)(123) <= estimated(414) xor estimated(415);
partial_sums(6)(124) <= estimated(94) xor estimated(95);
partial_sums(6)(125) <= estimated(350) xor estimated(351);
partial_sums(6)(126) <= estimated(222) xor estimated(223);
partial_sums(6)(127) <= estimated(478) xor estimated(479);
partial_sums(6)(128) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(129) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(130) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(131) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(132) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(133) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(134) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(135) <= estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(136) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(137) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(138) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(139) <= estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(140) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(141) <= estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(142) <= estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(143) <= estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(144) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(145) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(146) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(147) <= estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(148) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(149) <= estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(150) <= estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(151) <= estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(152) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(153) <= estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(154) <= estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(155) <= estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(156) <= estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(157) <= estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(158) <= estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(159) <= estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(160) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31);
partial_sums(6)(161) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287);
partial_sums(6)(162) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159);
partial_sums(6)(163) <= estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415);
partial_sums(6)(164) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95);
partial_sums(6)(165) <= estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351);
partial_sums(6)(166) <= estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223);
partial_sums(6)(167) <= estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479);
partial_sums(6)(168) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31);
partial_sums(6)(169) <= estimated(277) xor estimated(279) xor estimated(285) xor estimated(287);
partial_sums(6)(170) <= estimated(149) xor estimated(151) xor estimated(157) xor estimated(159);
partial_sums(6)(171) <= estimated(405) xor estimated(407) xor estimated(413) xor estimated(415);
partial_sums(6)(172) <= estimated(85) xor estimated(87) xor estimated(93) xor estimated(95);
partial_sums(6)(173) <= estimated(341) xor estimated(343) xor estimated(349) xor estimated(351);
partial_sums(6)(174) <= estimated(213) xor estimated(215) xor estimated(221) xor estimated(223);
partial_sums(6)(175) <= estimated(469) xor estimated(471) xor estimated(477) xor estimated(479);
partial_sums(6)(176) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31);
partial_sums(6)(177) <= estimated(269) xor estimated(271) xor estimated(285) xor estimated(287);
partial_sums(6)(178) <= estimated(141) xor estimated(143) xor estimated(157) xor estimated(159);
partial_sums(6)(179) <= estimated(397) xor estimated(399) xor estimated(413) xor estimated(415);
partial_sums(6)(180) <= estimated(77) xor estimated(79) xor estimated(93) xor estimated(95);
partial_sums(6)(181) <= estimated(333) xor estimated(335) xor estimated(349) xor estimated(351);
partial_sums(6)(182) <= estimated(205) xor estimated(207) xor estimated(221) xor estimated(223);
partial_sums(6)(183) <= estimated(461) xor estimated(463) xor estimated(477) xor estimated(479);
partial_sums(6)(184) <= estimated(29) xor estimated(31);
partial_sums(6)(185) <= estimated(285) xor estimated(287);
partial_sums(6)(186) <= estimated(157) xor estimated(159);
partial_sums(6)(187) <= estimated(413) xor estimated(415);
partial_sums(6)(188) <= estimated(93) xor estimated(95);
partial_sums(6)(189) <= estimated(349) xor estimated(351);
partial_sums(6)(190) <= estimated(221) xor estimated(223);
partial_sums(6)(191) <= estimated(477) xor estimated(479);
partial_sums(6)(192) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31);
partial_sums(6)(193) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287);
partial_sums(6)(194) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159);
partial_sums(6)(195) <= estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415);
partial_sums(6)(196) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95);
partial_sums(6)(197) <= estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351);
partial_sums(6)(198) <= estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223);
partial_sums(6)(199) <= estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479);
partial_sums(6)(200) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31);
partial_sums(6)(201) <= estimated(275) xor estimated(279) xor estimated(283) xor estimated(287);
partial_sums(6)(202) <= estimated(147) xor estimated(151) xor estimated(155) xor estimated(159);
partial_sums(6)(203) <= estimated(403) xor estimated(407) xor estimated(411) xor estimated(415);
partial_sums(6)(204) <= estimated(83) xor estimated(87) xor estimated(91) xor estimated(95);
partial_sums(6)(205) <= estimated(339) xor estimated(343) xor estimated(347) xor estimated(351);
partial_sums(6)(206) <= estimated(211) xor estimated(215) xor estimated(219) xor estimated(223);
partial_sums(6)(207) <= estimated(467) xor estimated(471) xor estimated(475) xor estimated(479);
partial_sums(6)(208) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31);
partial_sums(6)(209) <= estimated(267) xor estimated(271) xor estimated(283) xor estimated(287);
partial_sums(6)(210) <= estimated(139) xor estimated(143) xor estimated(155) xor estimated(159);
partial_sums(6)(211) <= estimated(395) xor estimated(399) xor estimated(411) xor estimated(415);
partial_sums(6)(212) <= estimated(75) xor estimated(79) xor estimated(91) xor estimated(95);
partial_sums(6)(213) <= estimated(331) xor estimated(335) xor estimated(347) xor estimated(351);
partial_sums(6)(214) <= estimated(203) xor estimated(207) xor estimated(219) xor estimated(223);
partial_sums(6)(215) <= estimated(459) xor estimated(463) xor estimated(475) xor estimated(479);
partial_sums(6)(216) <= estimated(27) xor estimated(31);
partial_sums(6)(217) <= estimated(283) xor estimated(287);
partial_sums(6)(218) <= estimated(155) xor estimated(159);
partial_sums(6)(219) <= estimated(411) xor estimated(415);
partial_sums(6)(220) <= estimated(91) xor estimated(95);
partial_sums(6)(221) <= estimated(347) xor estimated(351);
partial_sums(6)(222) <= estimated(219) xor estimated(223);
partial_sums(6)(223) <= estimated(475) xor estimated(479);
partial_sums(6)(224) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31);
partial_sums(6)(225) <= estimated(263) xor estimated(271) xor estimated(279) xor estimated(287);
partial_sums(6)(226) <= estimated(135) xor estimated(143) xor estimated(151) xor estimated(159);
partial_sums(6)(227) <= estimated(391) xor estimated(399) xor estimated(407) xor estimated(415);
partial_sums(6)(228) <= estimated(71) xor estimated(79) xor estimated(87) xor estimated(95);
partial_sums(6)(229) <= estimated(327) xor estimated(335) xor estimated(343) xor estimated(351);
partial_sums(6)(230) <= estimated(199) xor estimated(207) xor estimated(215) xor estimated(223);
partial_sums(6)(231) <= estimated(455) xor estimated(463) xor estimated(471) xor estimated(479);
partial_sums(6)(232) <= estimated(23) xor estimated(31);
partial_sums(6)(233) <= estimated(279) xor estimated(287);
partial_sums(6)(234) <= estimated(151) xor estimated(159);
partial_sums(6)(235) <= estimated(407) xor estimated(415);
partial_sums(6)(236) <= estimated(87) xor estimated(95);
partial_sums(6)(237) <= estimated(343) xor estimated(351);
partial_sums(6)(238) <= estimated(215) xor estimated(223);
partial_sums(6)(239) <= estimated(471) xor estimated(479);
partial_sums(6)(240) <= estimated(15) xor estimated(31);
partial_sums(6)(241) <= estimated(271) xor estimated(287);
partial_sums(6)(242) <= estimated(143) xor estimated(159);
partial_sums(6)(243) <= estimated(399) xor estimated(415);
partial_sums(6)(244) <= estimated(79) xor estimated(95);
partial_sums(6)(245) <= estimated(335) xor estimated(351);
partial_sums(6)(246) <= estimated(207) xor estimated(223);
partial_sums(6)(247) <= estimated(463) xor estimated(479);
partial_sums(6)(248) <= estimated(31);
partial_sums(6)(249) <= estimated(287);
partial_sums(6)(250) <= estimated(159);
partial_sums(6)(251) <= estimated(415);
partial_sums(6)(252) <= estimated(95);
partial_sums(6)(253) <= estimated(351);
partial_sums(6)(254) <= estimated(223);
partial_sums(6)(255) <= estimated(479);
partial_sums(7)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(1) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(2) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(3) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(4) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(5) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(6) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(7) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(8) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(9) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(10) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(11) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(12) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(13) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(14) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(15) <= estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(16) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(17) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(18) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(19) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(20) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(21) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(22) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(23) <= estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(24) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(25) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(26) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(27) <= estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(28) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(29) <= estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(30) <= estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(31) <= estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(32) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(33) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(34) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(35) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(36) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(37) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(38) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(39) <= estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(40) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(41) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(42) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(43) <= estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(44) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(45) <= estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(46) <= estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(47) <= estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(48) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(49) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(50) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(51) <= estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(52) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(53) <= estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(54) <= estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(55) <= estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(56) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(57) <= estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(58) <= estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(59) <= estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(60) <= estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(61) <= estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(62) <= estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(63) <= estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(64) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(65) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(66) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(67) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(68) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(69) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(70) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(71) <= estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(72) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(73) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(74) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(75) <= estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(76) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(77) <= estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(78) <= estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(79) <= estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(80) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(81) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(82) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(83) <= estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(84) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(85) <= estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(86) <= estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(87) <= estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(88) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(89) <= estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(90) <= estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(91) <= estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(92) <= estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(93) <= estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(94) <= estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(95) <= estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(96) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(97) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(98) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(99) <= estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(100) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(101) <= estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(102) <= estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(103) <= estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(104) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(105) <= estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(106) <= estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(107) <= estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(108) <= estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(109) <= estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(110) <= estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(111) <= estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(112) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31) xor estimated(46) xor estimated(47) xor estimated(62) xor estimated(63);
partial_sums(7)(113) <= estimated(270) xor estimated(271) xor estimated(286) xor estimated(287) xor estimated(302) xor estimated(303) xor estimated(318) xor estimated(319);
partial_sums(7)(114) <= estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191);
partial_sums(7)(115) <= estimated(398) xor estimated(399) xor estimated(414) xor estimated(415) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447);
partial_sums(7)(116) <= estimated(46) xor estimated(47) xor estimated(62) xor estimated(63);
partial_sums(7)(117) <= estimated(302) xor estimated(303) xor estimated(318) xor estimated(319);
partial_sums(7)(118) <= estimated(174) xor estimated(175) xor estimated(190) xor estimated(191);
partial_sums(7)(119) <= estimated(430) xor estimated(431) xor estimated(446) xor estimated(447);
partial_sums(7)(120) <= estimated(30) xor estimated(31) xor estimated(62) xor estimated(63);
partial_sums(7)(121) <= estimated(286) xor estimated(287) xor estimated(318) xor estimated(319);
partial_sums(7)(122) <= estimated(158) xor estimated(159) xor estimated(190) xor estimated(191);
partial_sums(7)(123) <= estimated(414) xor estimated(415) xor estimated(446) xor estimated(447);
partial_sums(7)(124) <= estimated(62) xor estimated(63);
partial_sums(7)(125) <= estimated(318) xor estimated(319);
partial_sums(7)(126) <= estimated(190) xor estimated(191);
partial_sums(7)(127) <= estimated(446) xor estimated(447);
partial_sums(7)(128) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(129) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(130) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(131) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(132) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(133) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(134) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(135) <= estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(136) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(137) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(138) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(139) <= estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(140) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(141) <= estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(142) <= estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(143) <= estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(144) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(145) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(146) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(147) <= estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(148) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(149) <= estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(150) <= estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(151) <= estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(152) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(153) <= estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(154) <= estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(155) <= estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(156) <= estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(157) <= estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(158) <= estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(159) <= estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(160) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(161) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(162) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(163) <= estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(164) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(165) <= estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(166) <= estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(167) <= estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(168) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(169) <= estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(170) <= estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(171) <= estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(172) <= estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(173) <= estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(174) <= estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(175) <= estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(176) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31) xor estimated(45) xor estimated(47) xor estimated(61) xor estimated(63);
partial_sums(7)(177) <= estimated(269) xor estimated(271) xor estimated(285) xor estimated(287) xor estimated(301) xor estimated(303) xor estimated(317) xor estimated(319);
partial_sums(7)(178) <= estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191);
partial_sums(7)(179) <= estimated(397) xor estimated(399) xor estimated(413) xor estimated(415) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447);
partial_sums(7)(180) <= estimated(45) xor estimated(47) xor estimated(61) xor estimated(63);
partial_sums(7)(181) <= estimated(301) xor estimated(303) xor estimated(317) xor estimated(319);
partial_sums(7)(182) <= estimated(173) xor estimated(175) xor estimated(189) xor estimated(191);
partial_sums(7)(183) <= estimated(429) xor estimated(431) xor estimated(445) xor estimated(447);
partial_sums(7)(184) <= estimated(29) xor estimated(31) xor estimated(61) xor estimated(63);
partial_sums(7)(185) <= estimated(285) xor estimated(287) xor estimated(317) xor estimated(319);
partial_sums(7)(186) <= estimated(157) xor estimated(159) xor estimated(189) xor estimated(191);
partial_sums(7)(187) <= estimated(413) xor estimated(415) xor estimated(445) xor estimated(447);
partial_sums(7)(188) <= estimated(61) xor estimated(63);
partial_sums(7)(189) <= estimated(317) xor estimated(319);
partial_sums(7)(190) <= estimated(189) xor estimated(191);
partial_sums(7)(191) <= estimated(445) xor estimated(447);
partial_sums(7)(192) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(193) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(194) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(195) <= estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(196) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(197) <= estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(198) <= estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(199) <= estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(200) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(201) <= estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(202) <= estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(203) <= estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(204) <= estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(205) <= estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(206) <= estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(207) <= estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(208) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31) xor estimated(43) xor estimated(47) xor estimated(59) xor estimated(63);
partial_sums(7)(209) <= estimated(267) xor estimated(271) xor estimated(283) xor estimated(287) xor estimated(299) xor estimated(303) xor estimated(315) xor estimated(319);
partial_sums(7)(210) <= estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191);
partial_sums(7)(211) <= estimated(395) xor estimated(399) xor estimated(411) xor estimated(415) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447);
partial_sums(7)(212) <= estimated(43) xor estimated(47) xor estimated(59) xor estimated(63);
partial_sums(7)(213) <= estimated(299) xor estimated(303) xor estimated(315) xor estimated(319);
partial_sums(7)(214) <= estimated(171) xor estimated(175) xor estimated(187) xor estimated(191);
partial_sums(7)(215) <= estimated(427) xor estimated(431) xor estimated(443) xor estimated(447);
partial_sums(7)(216) <= estimated(27) xor estimated(31) xor estimated(59) xor estimated(63);
partial_sums(7)(217) <= estimated(283) xor estimated(287) xor estimated(315) xor estimated(319);
partial_sums(7)(218) <= estimated(155) xor estimated(159) xor estimated(187) xor estimated(191);
partial_sums(7)(219) <= estimated(411) xor estimated(415) xor estimated(443) xor estimated(447);
partial_sums(7)(220) <= estimated(59) xor estimated(63);
partial_sums(7)(221) <= estimated(315) xor estimated(319);
partial_sums(7)(222) <= estimated(187) xor estimated(191);
partial_sums(7)(223) <= estimated(443) xor estimated(447);
partial_sums(7)(224) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31) xor estimated(39) xor estimated(47) xor estimated(55) xor estimated(63);
partial_sums(7)(225) <= estimated(263) xor estimated(271) xor estimated(279) xor estimated(287) xor estimated(295) xor estimated(303) xor estimated(311) xor estimated(319);
partial_sums(7)(226) <= estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191);
partial_sums(7)(227) <= estimated(391) xor estimated(399) xor estimated(407) xor estimated(415) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447);
partial_sums(7)(228) <= estimated(39) xor estimated(47) xor estimated(55) xor estimated(63);
partial_sums(7)(229) <= estimated(295) xor estimated(303) xor estimated(311) xor estimated(319);
partial_sums(7)(230) <= estimated(167) xor estimated(175) xor estimated(183) xor estimated(191);
partial_sums(7)(231) <= estimated(423) xor estimated(431) xor estimated(439) xor estimated(447);
partial_sums(7)(232) <= estimated(23) xor estimated(31) xor estimated(55) xor estimated(63);
partial_sums(7)(233) <= estimated(279) xor estimated(287) xor estimated(311) xor estimated(319);
partial_sums(7)(234) <= estimated(151) xor estimated(159) xor estimated(183) xor estimated(191);
partial_sums(7)(235) <= estimated(407) xor estimated(415) xor estimated(439) xor estimated(447);
partial_sums(7)(236) <= estimated(55) xor estimated(63);
partial_sums(7)(237) <= estimated(311) xor estimated(319);
partial_sums(7)(238) <= estimated(183) xor estimated(191);
partial_sums(7)(239) <= estimated(439) xor estimated(447);
partial_sums(7)(240) <= estimated(15) xor estimated(31) xor estimated(47) xor estimated(63);
partial_sums(7)(241) <= estimated(271) xor estimated(287) xor estimated(303) xor estimated(319);
partial_sums(7)(242) <= estimated(143) xor estimated(159) xor estimated(175) xor estimated(191);
partial_sums(7)(243) <= estimated(399) xor estimated(415) xor estimated(431) xor estimated(447);
partial_sums(7)(244) <= estimated(47) xor estimated(63);
partial_sums(7)(245) <= estimated(303) xor estimated(319);
partial_sums(7)(246) <= estimated(175) xor estimated(191);
partial_sums(7)(247) <= estimated(431) xor estimated(447);
partial_sums(7)(248) <= estimated(31) xor estimated(63);
partial_sums(7)(249) <= estimated(287) xor estimated(319);
partial_sums(7)(250) <= estimated(159) xor estimated(191);
partial_sums(7)(251) <= estimated(415) xor estimated(447);
partial_sums(7)(252) <= estimated(63);
partial_sums(7)(253) <= estimated(319);
partial_sums(7)(254) <= estimated(191);
partial_sums(7)(255) <= estimated(447);
partial_sums(8)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(1) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(2) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(3) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(4) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(5) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(6) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(7) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(8) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(9) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(10) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(11) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(12) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(13) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(14) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(15) <= estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(16) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(17) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(18) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(19) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(20) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(21) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(22) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(23) <= estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(24) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(25) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(26) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(27) <= estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(28) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(29) <= estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(30) <= estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(31) <= estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(32) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(33) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(34) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(35) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(36) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(37) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(38) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(39) <= estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(40) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(41) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(42) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(43) <= estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(44) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(45) <= estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(46) <= estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(47) <= estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(48) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(49) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(50) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(51) <= estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(52) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(53) <= estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(54) <= estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(55) <= estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(56) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(57) <= estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(58) <= estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(59) <= estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(60) <= estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(61) <= estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(62) <= estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(63) <= estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(64) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(65) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(66) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(67) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(68) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(69) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(70) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(71) <= estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(72) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(73) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(74) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(75) <= estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(76) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(77) <= estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(78) <= estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(79) <= estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(80) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(81) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(82) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(83) <= estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(84) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(85) <= estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(86) <= estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(87) <= estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(88) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(89) <= estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(90) <= estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(91) <= estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(92) <= estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(93) <= estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(94) <= estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(95) <= estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(96) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(97) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(98) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(99) <= estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(100) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(101) <= estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(102) <= estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(103) <= estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(104) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(105) <= estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(106) <= estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(107) <= estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(108) <= estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(109) <= estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(110) <= estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(111) <= estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(112) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31) xor estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(113) <= estimated(270) xor estimated(271) xor estimated(286) xor estimated(287) xor estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(114) <= estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(115) <= estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(116) <= estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(117) <= estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(118) <= estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(119) <= estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(120) <= estimated(30) xor estimated(31) xor estimated(62) xor estimated(63) xor estimated(94) xor estimated(95) xor estimated(126) xor estimated(127);
partial_sums(8)(121) <= estimated(286) xor estimated(287) xor estimated(318) xor estimated(319) xor estimated(350) xor estimated(351) xor estimated(382) xor estimated(383);
partial_sums(8)(122) <= estimated(94) xor estimated(95) xor estimated(126) xor estimated(127);
partial_sums(8)(123) <= estimated(350) xor estimated(351) xor estimated(382) xor estimated(383);
partial_sums(8)(124) <= estimated(62) xor estimated(63) xor estimated(126) xor estimated(127);
partial_sums(8)(125) <= estimated(318) xor estimated(319) xor estimated(382) xor estimated(383);
partial_sums(8)(126) <= estimated(126) xor estimated(127);
partial_sums(8)(127) <= estimated(382) xor estimated(383);
partial_sums(8)(128) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(129) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(130) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(131) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(132) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(133) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(134) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(135) <= estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(136) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(137) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(138) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(139) <= estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(140) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(141) <= estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(142) <= estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(143) <= estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(144) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(145) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(146) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(147) <= estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(148) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(149) <= estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(150) <= estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(151) <= estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(152) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(153) <= estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(154) <= estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(155) <= estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(156) <= estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(157) <= estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(158) <= estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(159) <= estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(160) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(161) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(162) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(163) <= estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(164) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(165) <= estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(166) <= estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(167) <= estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(168) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(169) <= estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(170) <= estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(171) <= estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(172) <= estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(173) <= estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(174) <= estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(175) <= estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(176) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31) xor estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(177) <= estimated(269) xor estimated(271) xor estimated(285) xor estimated(287) xor estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(178) <= estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(179) <= estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(180) <= estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(181) <= estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(182) <= estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(183) <= estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(184) <= estimated(29) xor estimated(31) xor estimated(61) xor estimated(63) xor estimated(93) xor estimated(95) xor estimated(125) xor estimated(127);
partial_sums(8)(185) <= estimated(285) xor estimated(287) xor estimated(317) xor estimated(319) xor estimated(349) xor estimated(351) xor estimated(381) xor estimated(383);
partial_sums(8)(186) <= estimated(93) xor estimated(95) xor estimated(125) xor estimated(127);
partial_sums(8)(187) <= estimated(349) xor estimated(351) xor estimated(381) xor estimated(383);
partial_sums(8)(188) <= estimated(61) xor estimated(63) xor estimated(125) xor estimated(127);
partial_sums(8)(189) <= estimated(317) xor estimated(319) xor estimated(381) xor estimated(383);
partial_sums(8)(190) <= estimated(125) xor estimated(127);
partial_sums(8)(191) <= estimated(381) xor estimated(383);
partial_sums(8)(192) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(193) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(194) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(195) <= estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(196) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(197) <= estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(198) <= estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(199) <= estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(200) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(201) <= estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(202) <= estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(203) <= estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(204) <= estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(205) <= estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(206) <= estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(207) <= estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(208) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31) xor estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(209) <= estimated(267) xor estimated(271) xor estimated(283) xor estimated(287) xor estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(210) <= estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(211) <= estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(212) <= estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(213) <= estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(214) <= estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(215) <= estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(216) <= estimated(27) xor estimated(31) xor estimated(59) xor estimated(63) xor estimated(91) xor estimated(95) xor estimated(123) xor estimated(127);
partial_sums(8)(217) <= estimated(283) xor estimated(287) xor estimated(315) xor estimated(319) xor estimated(347) xor estimated(351) xor estimated(379) xor estimated(383);
partial_sums(8)(218) <= estimated(91) xor estimated(95) xor estimated(123) xor estimated(127);
partial_sums(8)(219) <= estimated(347) xor estimated(351) xor estimated(379) xor estimated(383);
partial_sums(8)(220) <= estimated(59) xor estimated(63) xor estimated(123) xor estimated(127);
partial_sums(8)(221) <= estimated(315) xor estimated(319) xor estimated(379) xor estimated(383);
partial_sums(8)(222) <= estimated(123) xor estimated(127);
partial_sums(8)(223) <= estimated(379) xor estimated(383);
partial_sums(8)(224) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31) xor estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(225) <= estimated(263) xor estimated(271) xor estimated(279) xor estimated(287) xor estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(226) <= estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(227) <= estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(228) <= estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(229) <= estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(230) <= estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(231) <= estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(232) <= estimated(23) xor estimated(31) xor estimated(55) xor estimated(63) xor estimated(87) xor estimated(95) xor estimated(119) xor estimated(127);
partial_sums(8)(233) <= estimated(279) xor estimated(287) xor estimated(311) xor estimated(319) xor estimated(343) xor estimated(351) xor estimated(375) xor estimated(383);
partial_sums(8)(234) <= estimated(87) xor estimated(95) xor estimated(119) xor estimated(127);
partial_sums(8)(235) <= estimated(343) xor estimated(351) xor estimated(375) xor estimated(383);
partial_sums(8)(236) <= estimated(55) xor estimated(63) xor estimated(119) xor estimated(127);
partial_sums(8)(237) <= estimated(311) xor estimated(319) xor estimated(375) xor estimated(383);
partial_sums(8)(238) <= estimated(119) xor estimated(127);
partial_sums(8)(239) <= estimated(375) xor estimated(383);
partial_sums(8)(240) <= estimated(15) xor estimated(31) xor estimated(47) xor estimated(63) xor estimated(79) xor estimated(95) xor estimated(111) xor estimated(127);
partial_sums(8)(241) <= estimated(271) xor estimated(287) xor estimated(303) xor estimated(319) xor estimated(335) xor estimated(351) xor estimated(367) xor estimated(383);
partial_sums(8)(242) <= estimated(79) xor estimated(95) xor estimated(111) xor estimated(127);
partial_sums(8)(243) <= estimated(335) xor estimated(351) xor estimated(367) xor estimated(383);
partial_sums(8)(244) <= estimated(47) xor estimated(63) xor estimated(111) xor estimated(127);
partial_sums(8)(245) <= estimated(303) xor estimated(319) xor estimated(367) xor estimated(383);
partial_sums(8)(246) <= estimated(111) xor estimated(127);
partial_sums(8)(247) <= estimated(367) xor estimated(383);
partial_sums(8)(248) <= estimated(31) xor estimated(63) xor estimated(95) xor estimated(127);
partial_sums(8)(249) <= estimated(287) xor estimated(319) xor estimated(351) xor estimated(383);
partial_sums(8)(250) <= estimated(95) xor estimated(127);
partial_sums(8)(251) <= estimated(351) xor estimated(383);
partial_sums(8)(252) <= estimated(63) xor estimated(127);
partial_sums(8)(253) <= estimated(319) xor estimated(383);
partial_sums(8)(254) <= estimated(127);
partial_sums(8)(255) <= estimated(383);
partial_sums(9)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(1) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(2) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(3) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(4) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(5) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(6) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(7) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(8) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(9) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(10) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(11) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(12) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(13) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(14) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(15) <= estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(16) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(17) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(18) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(19) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(20) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(21) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(22) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(23) <= estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(24) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(25) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(26) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(27) <= estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(28) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(29) <= estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(30) <= estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(31) <= estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(32) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(33) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(34) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(35) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(36) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(37) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(38) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(39) <= estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(40) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(41) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(42) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(43) <= estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(44) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(45) <= estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(46) <= estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(47) <= estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(48) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(49) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(50) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(51) <= estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(52) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(53) <= estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(54) <= estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(55) <= estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(56) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(57) <= estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(58) <= estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(59) <= estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(60) <= estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(61) <= estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(62) <= estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(63) <= estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(64) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(65) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(66) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(67) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(68) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(69) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(70) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(71) <= estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(72) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(73) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(74) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(75) <= estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(76) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(77) <= estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(78) <= estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(79) <= estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(80) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(81) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(82) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(83) <= estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(84) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(85) <= estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(86) <= estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(87) <= estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(88) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(89) <= estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(90) <= estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(91) <= estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(92) <= estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(93) <= estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(94) <= estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(95) <= estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(96) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(97) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(98) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(99) <= estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(100) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(101) <= estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(102) <= estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(103) <= estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(104) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(105) <= estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(106) <= estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(107) <= estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(108) <= estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(109) <= estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(110) <= estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(111) <= estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(112) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31) xor estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(113) <= estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(114) <= estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(115) <= estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(116) <= estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(117) <= estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(118) <= estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(119) <= estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(120) <= estimated(30) xor estimated(31) xor estimated(62) xor estimated(63) xor estimated(94) xor estimated(95) xor estimated(126) xor estimated(127) xor estimated(158) xor estimated(159) xor estimated(190) xor estimated(191) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(121) <= estimated(158) xor estimated(159) xor estimated(190) xor estimated(191) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(122) <= estimated(94) xor estimated(95) xor estimated(126) xor estimated(127) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(123) <= estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(124) <= estimated(62) xor estimated(63) xor estimated(126) xor estimated(127) xor estimated(190) xor estimated(191) xor estimated(254) xor estimated(255);
partial_sums(9)(125) <= estimated(190) xor estimated(191) xor estimated(254) xor estimated(255);
partial_sums(9)(126) <= estimated(126) xor estimated(127) xor estimated(254) xor estimated(255);
partial_sums(9)(127) <= estimated(254) xor estimated(255);
partial_sums(9)(128) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(129) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(130) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(131) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(132) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(133) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(134) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(135) <= estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(136) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(137) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(138) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(139) <= estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(140) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(141) <= estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(142) <= estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(143) <= estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(144) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(145) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(146) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(147) <= estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(148) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(149) <= estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(150) <= estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(151) <= estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(152) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(153) <= estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(154) <= estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(155) <= estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(156) <= estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(157) <= estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(158) <= estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(159) <= estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(160) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(161) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(162) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(163) <= estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(164) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(165) <= estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(166) <= estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(167) <= estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(168) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(169) <= estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(170) <= estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(171) <= estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(172) <= estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(173) <= estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(174) <= estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(175) <= estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(176) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31) xor estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(177) <= estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(178) <= estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(179) <= estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(180) <= estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(181) <= estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(182) <= estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(183) <= estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(184) <= estimated(29) xor estimated(31) xor estimated(61) xor estimated(63) xor estimated(93) xor estimated(95) xor estimated(125) xor estimated(127) xor estimated(157) xor estimated(159) xor estimated(189) xor estimated(191) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(185) <= estimated(157) xor estimated(159) xor estimated(189) xor estimated(191) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(186) <= estimated(93) xor estimated(95) xor estimated(125) xor estimated(127) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(187) <= estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(188) <= estimated(61) xor estimated(63) xor estimated(125) xor estimated(127) xor estimated(189) xor estimated(191) xor estimated(253) xor estimated(255);
partial_sums(9)(189) <= estimated(189) xor estimated(191) xor estimated(253) xor estimated(255);
partial_sums(9)(190) <= estimated(125) xor estimated(127) xor estimated(253) xor estimated(255);
partial_sums(9)(191) <= estimated(253) xor estimated(255);
partial_sums(9)(192) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(193) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(194) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(195) <= estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(196) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(197) <= estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(198) <= estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(199) <= estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(200) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(201) <= estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(202) <= estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(203) <= estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(204) <= estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(205) <= estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(206) <= estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(207) <= estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(208) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31) xor estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(209) <= estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(210) <= estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(211) <= estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(212) <= estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(213) <= estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(214) <= estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(215) <= estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(216) <= estimated(27) xor estimated(31) xor estimated(59) xor estimated(63) xor estimated(91) xor estimated(95) xor estimated(123) xor estimated(127) xor estimated(155) xor estimated(159) xor estimated(187) xor estimated(191) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(217) <= estimated(155) xor estimated(159) xor estimated(187) xor estimated(191) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(218) <= estimated(91) xor estimated(95) xor estimated(123) xor estimated(127) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(219) <= estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(220) <= estimated(59) xor estimated(63) xor estimated(123) xor estimated(127) xor estimated(187) xor estimated(191) xor estimated(251) xor estimated(255);
partial_sums(9)(221) <= estimated(187) xor estimated(191) xor estimated(251) xor estimated(255);
partial_sums(9)(222) <= estimated(123) xor estimated(127) xor estimated(251) xor estimated(255);
partial_sums(9)(223) <= estimated(251) xor estimated(255);
partial_sums(9)(224) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31) xor estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(225) <= estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(226) <= estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(227) <= estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(228) <= estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(229) <= estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(230) <= estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(231) <= estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(232) <= estimated(23) xor estimated(31) xor estimated(55) xor estimated(63) xor estimated(87) xor estimated(95) xor estimated(119) xor estimated(127) xor estimated(151) xor estimated(159) xor estimated(183) xor estimated(191) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(233) <= estimated(151) xor estimated(159) xor estimated(183) xor estimated(191) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(234) <= estimated(87) xor estimated(95) xor estimated(119) xor estimated(127) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(235) <= estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(236) <= estimated(55) xor estimated(63) xor estimated(119) xor estimated(127) xor estimated(183) xor estimated(191) xor estimated(247) xor estimated(255);
partial_sums(9)(237) <= estimated(183) xor estimated(191) xor estimated(247) xor estimated(255);
partial_sums(9)(238) <= estimated(119) xor estimated(127) xor estimated(247) xor estimated(255);
partial_sums(9)(239) <= estimated(247) xor estimated(255);
partial_sums(9)(240) <= estimated(15) xor estimated(31) xor estimated(47) xor estimated(63) xor estimated(79) xor estimated(95) xor estimated(111) xor estimated(127) xor estimated(143) xor estimated(159) xor estimated(175) xor estimated(191) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(241) <= estimated(143) xor estimated(159) xor estimated(175) xor estimated(191) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(242) <= estimated(79) xor estimated(95) xor estimated(111) xor estimated(127) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(243) <= estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(244) <= estimated(47) xor estimated(63) xor estimated(111) xor estimated(127) xor estimated(175) xor estimated(191) xor estimated(239) xor estimated(255);
partial_sums(9)(245) <= estimated(175) xor estimated(191) xor estimated(239) xor estimated(255);
partial_sums(9)(246) <= estimated(111) xor estimated(127) xor estimated(239) xor estimated(255);
partial_sums(9)(247) <= estimated(239) xor estimated(255);
partial_sums(9)(248) <= estimated(31) xor estimated(63) xor estimated(95) xor estimated(127) xor estimated(159) xor estimated(191) xor estimated(223) xor estimated(255);
partial_sums(9)(249) <= estimated(159) xor estimated(191) xor estimated(223) xor estimated(255);
partial_sums(9)(250) <= estimated(95) xor estimated(127) xor estimated(223) xor estimated(255);
partial_sums(9)(251) <= estimated(223) xor estimated(255);
partial_sums(9)(252) <= estimated(63) xor estimated(127) xor estimated(191) xor estimated(255);
partial_sums(9)(253) <= estimated(191) xor estimated(255);
partial_sums(9)(254) <= estimated(127) xor estimated(255);
partial_sums(9)(255) <= estimated(255);
end Behavioral;


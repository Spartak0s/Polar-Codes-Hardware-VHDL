----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:50:12 04/01/2016 
-- Design Name: 
-- Module Name:    Decoder1024 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.all;
use work.MyPackage.all;
use IEEE.math_real.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Decoder1024 is
    Port ( clk : in  STD_LOGIC;
			  rst: in STD_LOGIC;
			  ce_inputs: in STD_LOGIC;
			  inputs : in data;
           outputs : out  STD_LOGIC_VECTOR (N/2-1 downto 0));
end Decoder1024;

architecture Behavioral of Decoder1024 is
	signal P: llr_2d := (others=>(others=>(others=> '0')));
	signal u : std_logic_vector(N-2 downto 0) := (others => '0');
	signal s: s_2d := (others=>(others=> '0'));
	signal ce_outputs : std_logic := '1';
begin
	--Input Registers
	GEN_REG_INPUT:
	for I in 0 to N-1 generate
		U_D_FF_Inputs: entity work.D_FF_gen generic map(width=>integer_part+fractional_part)
										 port map(clk =>clk,
													 rst =>rst,
													 ce =>ce_inputs,
													 d =>inputs(I),
													 q =>P(stages)(I));
	end generate GEN_REG_INPUT;
	
--	GEN_STAGES:
--	
--	for I in 1 to stages-1 generate
--		for J in 0 to 1023 generate
--			if (((J / MOD(2**(I-1),2))) == 0)
--				F: entity work.F port map(P(I)(J)
--		end generate;
--	end generate;
-- STAGE 9
U_F100: entity F port map(lamdaA => P(10)(0),lamdaB => P(10)(1),lamdaOut => P(9)(0));
U_G101: entity G port map(lamdaA => P(10)(0),lamdaB => P(10)(1),s => s(10)(0),lamdaOut => P(9)(1));
U_F102: entity F port map(lamdaA => P(10)(2),lamdaB => P(10)(3),lamdaOut => P(9)(2));
U_G103: entity G port map(lamdaA => P(10)(2),lamdaB => P(10)(3),s => s(10)(1),lamdaOut => P(9)(3));
U_F104: entity F port map(lamdaA => P(10)(4),lamdaB => P(10)(5),lamdaOut => P(9)(4));
U_G105: entity G port map(lamdaA => P(10)(4),lamdaB => P(10)(5),s => s(10)(2),lamdaOut => P(9)(5));
U_F106: entity F port map(lamdaA => P(10)(6),lamdaB => P(10)(7),lamdaOut => P(9)(6));
U_G107: entity G port map(lamdaA => P(10)(6),lamdaB => P(10)(7),s => s(10)(3),lamdaOut => P(9)(7));
U_F108: entity F port map(lamdaA => P(10)(8),lamdaB => P(10)(9),lamdaOut => P(9)(8));
U_G109: entity G port map(lamdaA => P(10)(8),lamdaB => P(10)(9),s => s(10)(4),lamdaOut => P(9)(9));
U_F1010: entity F port map(lamdaA => P(10)(10),lamdaB => P(10)(11),lamdaOut => P(9)(10));
U_G1011: entity G port map(lamdaA => P(10)(10),lamdaB => P(10)(11),s => s(10)(5),lamdaOut => P(9)(11));
U_F1012: entity F port map(lamdaA => P(10)(12),lamdaB => P(10)(13),lamdaOut => P(9)(12));
U_G1013: entity G port map(lamdaA => P(10)(12),lamdaB => P(10)(13),s => s(10)(6),lamdaOut => P(9)(13));
U_F1014: entity F port map(lamdaA => P(10)(14),lamdaB => P(10)(15),lamdaOut => P(9)(14));
U_G1015: entity G port map(lamdaA => P(10)(14),lamdaB => P(10)(15),s => s(10)(7),lamdaOut => P(9)(15));
U_F1016: entity F port map(lamdaA => P(10)(16),lamdaB => P(10)(17),lamdaOut => P(9)(16));
U_G1017: entity G port map(lamdaA => P(10)(16),lamdaB => P(10)(17),s => s(10)(8),lamdaOut => P(9)(17));
U_F1018: entity F port map(lamdaA => P(10)(18),lamdaB => P(10)(19),lamdaOut => P(9)(18));
U_G1019: entity G port map(lamdaA => P(10)(18),lamdaB => P(10)(19),s => s(10)(9),lamdaOut => P(9)(19));
U_F1020: entity F port map(lamdaA => P(10)(20),lamdaB => P(10)(21),lamdaOut => P(9)(20));
U_G1021: entity G port map(lamdaA => P(10)(20),lamdaB => P(10)(21),s => s(10)(10),lamdaOut => P(9)(21));
U_F1022: entity F port map(lamdaA => P(10)(22),lamdaB => P(10)(23),lamdaOut => P(9)(22));
U_G1023: entity G port map(lamdaA => P(10)(22),lamdaB => P(10)(23),s => s(10)(11),lamdaOut => P(9)(23));
U_F1024: entity F port map(lamdaA => P(10)(24),lamdaB => P(10)(25),lamdaOut => P(9)(24));
U_G1025: entity G port map(lamdaA => P(10)(24),lamdaB => P(10)(25),s => s(10)(12),lamdaOut => P(9)(25));
U_F1026: entity F port map(lamdaA => P(10)(26),lamdaB => P(10)(27),lamdaOut => P(9)(26));
U_G1027: entity G port map(lamdaA => P(10)(26),lamdaB => P(10)(27),s => s(10)(13),lamdaOut => P(9)(27));
U_F1028: entity F port map(lamdaA => P(10)(28),lamdaB => P(10)(29),lamdaOut => P(9)(28));
U_G1029: entity G port map(lamdaA => P(10)(28),lamdaB => P(10)(29),s => s(10)(14),lamdaOut => P(9)(29));
U_F1030: entity F port map(lamdaA => P(10)(30),lamdaB => P(10)(31),lamdaOut => P(9)(30));
U_G1031: entity G port map(lamdaA => P(10)(30),lamdaB => P(10)(31),s => s(10)(15),lamdaOut => P(9)(31));
U_F1032: entity F port map(lamdaA => P(10)(32),lamdaB => P(10)(33),lamdaOut => P(9)(32));
U_G1033: entity G port map(lamdaA => P(10)(32),lamdaB => P(10)(33),s => s(10)(16),lamdaOut => P(9)(33));
U_F1034: entity F port map(lamdaA => P(10)(34),lamdaB => P(10)(35),lamdaOut => P(9)(34));
U_G1035: entity G port map(lamdaA => P(10)(34),lamdaB => P(10)(35),s => s(10)(17),lamdaOut => P(9)(35));
U_F1036: entity F port map(lamdaA => P(10)(36),lamdaB => P(10)(37),lamdaOut => P(9)(36));
U_G1037: entity G port map(lamdaA => P(10)(36),lamdaB => P(10)(37),s => s(10)(18),lamdaOut => P(9)(37));
U_F1038: entity F port map(lamdaA => P(10)(38),lamdaB => P(10)(39),lamdaOut => P(9)(38));
U_G1039: entity G port map(lamdaA => P(10)(38),lamdaB => P(10)(39),s => s(10)(19),lamdaOut => P(9)(39));
U_F1040: entity F port map(lamdaA => P(10)(40),lamdaB => P(10)(41),lamdaOut => P(9)(40));
U_G1041: entity G port map(lamdaA => P(10)(40),lamdaB => P(10)(41),s => s(10)(20),lamdaOut => P(9)(41));
U_F1042: entity F port map(lamdaA => P(10)(42),lamdaB => P(10)(43),lamdaOut => P(9)(42));
U_G1043: entity G port map(lamdaA => P(10)(42),lamdaB => P(10)(43),s => s(10)(21),lamdaOut => P(9)(43));
U_F1044: entity F port map(lamdaA => P(10)(44),lamdaB => P(10)(45),lamdaOut => P(9)(44));
U_G1045: entity G port map(lamdaA => P(10)(44),lamdaB => P(10)(45),s => s(10)(22),lamdaOut => P(9)(45));
U_F1046: entity F port map(lamdaA => P(10)(46),lamdaB => P(10)(47),lamdaOut => P(9)(46));
U_G1047: entity G port map(lamdaA => P(10)(46),lamdaB => P(10)(47),s => s(10)(23),lamdaOut => P(9)(47));
U_F1048: entity F port map(lamdaA => P(10)(48),lamdaB => P(10)(49),lamdaOut => P(9)(48));
U_G1049: entity G port map(lamdaA => P(10)(48),lamdaB => P(10)(49),s => s(10)(24),lamdaOut => P(9)(49));
U_F1050: entity F port map(lamdaA => P(10)(50),lamdaB => P(10)(51),lamdaOut => P(9)(50));
U_G1051: entity G port map(lamdaA => P(10)(50),lamdaB => P(10)(51),s => s(10)(25),lamdaOut => P(9)(51));
U_F1052: entity F port map(lamdaA => P(10)(52),lamdaB => P(10)(53),lamdaOut => P(9)(52));
U_G1053: entity G port map(lamdaA => P(10)(52),lamdaB => P(10)(53),s => s(10)(26),lamdaOut => P(9)(53));
U_F1054: entity F port map(lamdaA => P(10)(54),lamdaB => P(10)(55),lamdaOut => P(9)(54));
U_G1055: entity G port map(lamdaA => P(10)(54),lamdaB => P(10)(55),s => s(10)(27),lamdaOut => P(9)(55));
U_F1056: entity F port map(lamdaA => P(10)(56),lamdaB => P(10)(57),lamdaOut => P(9)(56));
U_G1057: entity G port map(lamdaA => P(10)(56),lamdaB => P(10)(57),s => s(10)(28),lamdaOut => P(9)(57));
U_F1058: entity F port map(lamdaA => P(10)(58),lamdaB => P(10)(59),lamdaOut => P(9)(58));
U_G1059: entity G port map(lamdaA => P(10)(58),lamdaB => P(10)(59),s => s(10)(29),lamdaOut => P(9)(59));
U_F1060: entity F port map(lamdaA => P(10)(60),lamdaB => P(10)(61),lamdaOut => P(9)(60));
U_G1061: entity G port map(lamdaA => P(10)(60),lamdaB => P(10)(61),s => s(10)(30),lamdaOut => P(9)(61));
U_F1062: entity F port map(lamdaA => P(10)(62),lamdaB => P(10)(63),lamdaOut => P(9)(62));
U_G1063: entity G port map(lamdaA => P(10)(62),lamdaB => P(10)(63),s => s(10)(31),lamdaOut => P(9)(63));
U_F1064: entity F port map(lamdaA => P(10)(64),lamdaB => P(10)(65),lamdaOut => P(9)(64));
U_G1065: entity G port map(lamdaA => P(10)(64),lamdaB => P(10)(65),s => s(10)(32),lamdaOut => P(9)(65));
U_F1066: entity F port map(lamdaA => P(10)(66),lamdaB => P(10)(67),lamdaOut => P(9)(66));
U_G1067: entity G port map(lamdaA => P(10)(66),lamdaB => P(10)(67),s => s(10)(33),lamdaOut => P(9)(67));
U_F1068: entity F port map(lamdaA => P(10)(68),lamdaB => P(10)(69),lamdaOut => P(9)(68));
U_G1069: entity G port map(lamdaA => P(10)(68),lamdaB => P(10)(69),s => s(10)(34),lamdaOut => P(9)(69));
U_F1070: entity F port map(lamdaA => P(10)(70),lamdaB => P(10)(71),lamdaOut => P(9)(70));
U_G1071: entity G port map(lamdaA => P(10)(70),lamdaB => P(10)(71),s => s(10)(35),lamdaOut => P(9)(71));
U_F1072: entity F port map(lamdaA => P(10)(72),lamdaB => P(10)(73),lamdaOut => P(9)(72));
U_G1073: entity G port map(lamdaA => P(10)(72),lamdaB => P(10)(73),s => s(10)(36),lamdaOut => P(9)(73));
U_F1074: entity F port map(lamdaA => P(10)(74),lamdaB => P(10)(75),lamdaOut => P(9)(74));
U_G1075: entity G port map(lamdaA => P(10)(74),lamdaB => P(10)(75),s => s(10)(37),lamdaOut => P(9)(75));
U_F1076: entity F port map(lamdaA => P(10)(76),lamdaB => P(10)(77),lamdaOut => P(9)(76));
U_G1077: entity G port map(lamdaA => P(10)(76),lamdaB => P(10)(77),s => s(10)(38),lamdaOut => P(9)(77));
U_F1078: entity F port map(lamdaA => P(10)(78),lamdaB => P(10)(79),lamdaOut => P(9)(78));
U_G1079: entity G port map(lamdaA => P(10)(78),lamdaB => P(10)(79),s => s(10)(39),lamdaOut => P(9)(79));
U_F1080: entity F port map(lamdaA => P(10)(80),lamdaB => P(10)(81),lamdaOut => P(9)(80));
U_G1081: entity G port map(lamdaA => P(10)(80),lamdaB => P(10)(81),s => s(10)(40),lamdaOut => P(9)(81));
U_F1082: entity F port map(lamdaA => P(10)(82),lamdaB => P(10)(83),lamdaOut => P(9)(82));
U_G1083: entity G port map(lamdaA => P(10)(82),lamdaB => P(10)(83),s => s(10)(41),lamdaOut => P(9)(83));
U_F1084: entity F port map(lamdaA => P(10)(84),lamdaB => P(10)(85),lamdaOut => P(9)(84));
U_G1085: entity G port map(lamdaA => P(10)(84),lamdaB => P(10)(85),s => s(10)(42),lamdaOut => P(9)(85));
U_F1086: entity F port map(lamdaA => P(10)(86),lamdaB => P(10)(87),lamdaOut => P(9)(86));
U_G1087: entity G port map(lamdaA => P(10)(86),lamdaB => P(10)(87),s => s(10)(43),lamdaOut => P(9)(87));
U_F1088: entity F port map(lamdaA => P(10)(88),lamdaB => P(10)(89),lamdaOut => P(9)(88));
U_G1089: entity G port map(lamdaA => P(10)(88),lamdaB => P(10)(89),s => s(10)(44),lamdaOut => P(9)(89));
U_F1090: entity F port map(lamdaA => P(10)(90),lamdaB => P(10)(91),lamdaOut => P(9)(90));
U_G1091: entity G port map(lamdaA => P(10)(90),lamdaB => P(10)(91),s => s(10)(45),lamdaOut => P(9)(91));
U_F1092: entity F port map(lamdaA => P(10)(92),lamdaB => P(10)(93),lamdaOut => P(9)(92));
U_G1093: entity G port map(lamdaA => P(10)(92),lamdaB => P(10)(93),s => s(10)(46),lamdaOut => P(9)(93));
U_F1094: entity F port map(lamdaA => P(10)(94),lamdaB => P(10)(95),lamdaOut => P(9)(94));
U_G1095: entity G port map(lamdaA => P(10)(94),lamdaB => P(10)(95),s => s(10)(47),lamdaOut => P(9)(95));
U_F1096: entity F port map(lamdaA => P(10)(96),lamdaB => P(10)(97),lamdaOut => P(9)(96));
U_G1097: entity G port map(lamdaA => P(10)(96),lamdaB => P(10)(97),s => s(10)(48),lamdaOut => P(9)(97));
U_F1098: entity F port map(lamdaA => P(10)(98),lamdaB => P(10)(99),lamdaOut => P(9)(98));
U_G1099: entity G port map(lamdaA => P(10)(98),lamdaB => P(10)(99),s => s(10)(49),lamdaOut => P(9)(99));
U_F10100: entity F port map(lamdaA => P(10)(100),lamdaB => P(10)(101),lamdaOut => P(9)(100));
U_G10101: entity G port map(lamdaA => P(10)(100),lamdaB => P(10)(101),s => s(10)(50),lamdaOut => P(9)(101));
U_F10102: entity F port map(lamdaA => P(10)(102),lamdaB => P(10)(103),lamdaOut => P(9)(102));
U_G10103: entity G port map(lamdaA => P(10)(102),lamdaB => P(10)(103),s => s(10)(51),lamdaOut => P(9)(103));
U_F10104: entity F port map(lamdaA => P(10)(104),lamdaB => P(10)(105),lamdaOut => P(9)(104));
U_G10105: entity G port map(lamdaA => P(10)(104),lamdaB => P(10)(105),s => s(10)(52),lamdaOut => P(9)(105));
U_F10106: entity F port map(lamdaA => P(10)(106),lamdaB => P(10)(107),lamdaOut => P(9)(106));
U_G10107: entity G port map(lamdaA => P(10)(106),lamdaB => P(10)(107),s => s(10)(53),lamdaOut => P(9)(107));
U_F10108: entity F port map(lamdaA => P(10)(108),lamdaB => P(10)(109),lamdaOut => P(9)(108));
U_G10109: entity G port map(lamdaA => P(10)(108),lamdaB => P(10)(109),s => s(10)(54),lamdaOut => P(9)(109));
U_F10110: entity F port map(lamdaA => P(10)(110),lamdaB => P(10)(111),lamdaOut => P(9)(110));
U_G10111: entity G port map(lamdaA => P(10)(110),lamdaB => P(10)(111),s => s(10)(55),lamdaOut => P(9)(111));
U_F10112: entity F port map(lamdaA => P(10)(112),lamdaB => P(10)(113),lamdaOut => P(9)(112));
U_G10113: entity G port map(lamdaA => P(10)(112),lamdaB => P(10)(113),s => s(10)(56),lamdaOut => P(9)(113));
U_F10114: entity F port map(lamdaA => P(10)(114),lamdaB => P(10)(115),lamdaOut => P(9)(114));
U_G10115: entity G port map(lamdaA => P(10)(114),lamdaB => P(10)(115),s => s(10)(57),lamdaOut => P(9)(115));
U_F10116: entity F port map(lamdaA => P(10)(116),lamdaB => P(10)(117),lamdaOut => P(9)(116));
U_G10117: entity G port map(lamdaA => P(10)(116),lamdaB => P(10)(117),s => s(10)(58),lamdaOut => P(9)(117));
U_F10118: entity F port map(lamdaA => P(10)(118),lamdaB => P(10)(119),lamdaOut => P(9)(118));
U_G10119: entity G port map(lamdaA => P(10)(118),lamdaB => P(10)(119),s => s(10)(59),lamdaOut => P(9)(119));
U_F10120: entity F port map(lamdaA => P(10)(120),lamdaB => P(10)(121),lamdaOut => P(9)(120));
U_G10121: entity G port map(lamdaA => P(10)(120),lamdaB => P(10)(121),s => s(10)(60),lamdaOut => P(9)(121));
U_F10122: entity F port map(lamdaA => P(10)(122),lamdaB => P(10)(123),lamdaOut => P(9)(122));
U_G10123: entity G port map(lamdaA => P(10)(122),lamdaB => P(10)(123),s => s(10)(61),lamdaOut => P(9)(123));
U_F10124: entity F port map(lamdaA => P(10)(124),lamdaB => P(10)(125),lamdaOut => P(9)(124));
U_G10125: entity G port map(lamdaA => P(10)(124),lamdaB => P(10)(125),s => s(10)(62),lamdaOut => P(9)(125));
U_F10126: entity F port map(lamdaA => P(10)(126),lamdaB => P(10)(127),lamdaOut => P(9)(126));
U_G10127: entity G port map(lamdaA => P(10)(126),lamdaB => P(10)(127),s => s(10)(63),lamdaOut => P(9)(127));
U_F10128: entity F port map(lamdaA => P(10)(128),lamdaB => P(10)(129),lamdaOut => P(9)(128));
U_G10129: entity G port map(lamdaA => P(10)(128),lamdaB => P(10)(129),s => s(10)(64),lamdaOut => P(9)(129));
U_F10130: entity F port map(lamdaA => P(10)(130),lamdaB => P(10)(131),lamdaOut => P(9)(130));
U_G10131: entity G port map(lamdaA => P(10)(130),lamdaB => P(10)(131),s => s(10)(65),lamdaOut => P(9)(131));
U_F10132: entity F port map(lamdaA => P(10)(132),lamdaB => P(10)(133),lamdaOut => P(9)(132));
U_G10133: entity G port map(lamdaA => P(10)(132),lamdaB => P(10)(133),s => s(10)(66),lamdaOut => P(9)(133));
U_F10134: entity F port map(lamdaA => P(10)(134),lamdaB => P(10)(135),lamdaOut => P(9)(134));
U_G10135: entity G port map(lamdaA => P(10)(134),lamdaB => P(10)(135),s => s(10)(67),lamdaOut => P(9)(135));
U_F10136: entity F port map(lamdaA => P(10)(136),lamdaB => P(10)(137),lamdaOut => P(9)(136));
U_G10137: entity G port map(lamdaA => P(10)(136),lamdaB => P(10)(137),s => s(10)(68),lamdaOut => P(9)(137));
U_F10138: entity F port map(lamdaA => P(10)(138),lamdaB => P(10)(139),lamdaOut => P(9)(138));
U_G10139: entity G port map(lamdaA => P(10)(138),lamdaB => P(10)(139),s => s(10)(69),lamdaOut => P(9)(139));
U_F10140: entity F port map(lamdaA => P(10)(140),lamdaB => P(10)(141),lamdaOut => P(9)(140));
U_G10141: entity G port map(lamdaA => P(10)(140),lamdaB => P(10)(141),s => s(10)(70),lamdaOut => P(9)(141));
U_F10142: entity F port map(lamdaA => P(10)(142),lamdaB => P(10)(143),lamdaOut => P(9)(142));
U_G10143: entity G port map(lamdaA => P(10)(142),lamdaB => P(10)(143),s => s(10)(71),lamdaOut => P(9)(143));
U_F10144: entity F port map(lamdaA => P(10)(144),lamdaB => P(10)(145),lamdaOut => P(9)(144));
U_G10145: entity G port map(lamdaA => P(10)(144),lamdaB => P(10)(145),s => s(10)(72),lamdaOut => P(9)(145));
U_F10146: entity F port map(lamdaA => P(10)(146),lamdaB => P(10)(147),lamdaOut => P(9)(146));
U_G10147: entity G port map(lamdaA => P(10)(146),lamdaB => P(10)(147),s => s(10)(73),lamdaOut => P(9)(147));
U_F10148: entity F port map(lamdaA => P(10)(148),lamdaB => P(10)(149),lamdaOut => P(9)(148));
U_G10149: entity G port map(lamdaA => P(10)(148),lamdaB => P(10)(149),s => s(10)(74),lamdaOut => P(9)(149));
U_F10150: entity F port map(lamdaA => P(10)(150),lamdaB => P(10)(151),lamdaOut => P(9)(150));
U_G10151: entity G port map(lamdaA => P(10)(150),lamdaB => P(10)(151),s => s(10)(75),lamdaOut => P(9)(151));
U_F10152: entity F port map(lamdaA => P(10)(152),lamdaB => P(10)(153),lamdaOut => P(9)(152));
U_G10153: entity G port map(lamdaA => P(10)(152),lamdaB => P(10)(153),s => s(10)(76),lamdaOut => P(9)(153));
U_F10154: entity F port map(lamdaA => P(10)(154),lamdaB => P(10)(155),lamdaOut => P(9)(154));
U_G10155: entity G port map(lamdaA => P(10)(154),lamdaB => P(10)(155),s => s(10)(77),lamdaOut => P(9)(155));
U_F10156: entity F port map(lamdaA => P(10)(156),lamdaB => P(10)(157),lamdaOut => P(9)(156));
U_G10157: entity G port map(lamdaA => P(10)(156),lamdaB => P(10)(157),s => s(10)(78),lamdaOut => P(9)(157));
U_F10158: entity F port map(lamdaA => P(10)(158),lamdaB => P(10)(159),lamdaOut => P(9)(158));
U_G10159: entity G port map(lamdaA => P(10)(158),lamdaB => P(10)(159),s => s(10)(79),lamdaOut => P(9)(159));
U_F10160: entity F port map(lamdaA => P(10)(160),lamdaB => P(10)(161),lamdaOut => P(9)(160));
U_G10161: entity G port map(lamdaA => P(10)(160),lamdaB => P(10)(161),s => s(10)(80),lamdaOut => P(9)(161));
U_F10162: entity F port map(lamdaA => P(10)(162),lamdaB => P(10)(163),lamdaOut => P(9)(162));
U_G10163: entity G port map(lamdaA => P(10)(162),lamdaB => P(10)(163),s => s(10)(81),lamdaOut => P(9)(163));
U_F10164: entity F port map(lamdaA => P(10)(164),lamdaB => P(10)(165),lamdaOut => P(9)(164));
U_G10165: entity G port map(lamdaA => P(10)(164),lamdaB => P(10)(165),s => s(10)(82),lamdaOut => P(9)(165));
U_F10166: entity F port map(lamdaA => P(10)(166),lamdaB => P(10)(167),lamdaOut => P(9)(166));
U_G10167: entity G port map(lamdaA => P(10)(166),lamdaB => P(10)(167),s => s(10)(83),lamdaOut => P(9)(167));
U_F10168: entity F port map(lamdaA => P(10)(168),lamdaB => P(10)(169),lamdaOut => P(9)(168));
U_G10169: entity G port map(lamdaA => P(10)(168),lamdaB => P(10)(169),s => s(10)(84),lamdaOut => P(9)(169));
U_F10170: entity F port map(lamdaA => P(10)(170),lamdaB => P(10)(171),lamdaOut => P(9)(170));
U_G10171: entity G port map(lamdaA => P(10)(170),lamdaB => P(10)(171),s => s(10)(85),lamdaOut => P(9)(171));
U_F10172: entity F port map(lamdaA => P(10)(172),lamdaB => P(10)(173),lamdaOut => P(9)(172));
U_G10173: entity G port map(lamdaA => P(10)(172),lamdaB => P(10)(173),s => s(10)(86),lamdaOut => P(9)(173));
U_F10174: entity F port map(lamdaA => P(10)(174),lamdaB => P(10)(175),lamdaOut => P(9)(174));
U_G10175: entity G port map(lamdaA => P(10)(174),lamdaB => P(10)(175),s => s(10)(87),lamdaOut => P(9)(175));
U_F10176: entity F port map(lamdaA => P(10)(176),lamdaB => P(10)(177),lamdaOut => P(9)(176));
U_G10177: entity G port map(lamdaA => P(10)(176),lamdaB => P(10)(177),s => s(10)(88),lamdaOut => P(9)(177));
U_F10178: entity F port map(lamdaA => P(10)(178),lamdaB => P(10)(179),lamdaOut => P(9)(178));
U_G10179: entity G port map(lamdaA => P(10)(178),lamdaB => P(10)(179),s => s(10)(89),lamdaOut => P(9)(179));
U_F10180: entity F port map(lamdaA => P(10)(180),lamdaB => P(10)(181),lamdaOut => P(9)(180));
U_G10181: entity G port map(lamdaA => P(10)(180),lamdaB => P(10)(181),s => s(10)(90),lamdaOut => P(9)(181));
U_F10182: entity F port map(lamdaA => P(10)(182),lamdaB => P(10)(183),lamdaOut => P(9)(182));
U_G10183: entity G port map(lamdaA => P(10)(182),lamdaB => P(10)(183),s => s(10)(91),lamdaOut => P(9)(183));
U_F10184: entity F port map(lamdaA => P(10)(184),lamdaB => P(10)(185),lamdaOut => P(9)(184));
U_G10185: entity G port map(lamdaA => P(10)(184),lamdaB => P(10)(185),s => s(10)(92),lamdaOut => P(9)(185));
U_F10186: entity F port map(lamdaA => P(10)(186),lamdaB => P(10)(187),lamdaOut => P(9)(186));
U_G10187: entity G port map(lamdaA => P(10)(186),lamdaB => P(10)(187),s => s(10)(93),lamdaOut => P(9)(187));
U_F10188: entity F port map(lamdaA => P(10)(188),lamdaB => P(10)(189),lamdaOut => P(9)(188));
U_G10189: entity G port map(lamdaA => P(10)(188),lamdaB => P(10)(189),s => s(10)(94),lamdaOut => P(9)(189));
U_F10190: entity F port map(lamdaA => P(10)(190),lamdaB => P(10)(191),lamdaOut => P(9)(190));
U_G10191: entity G port map(lamdaA => P(10)(190),lamdaB => P(10)(191),s => s(10)(95),lamdaOut => P(9)(191));
U_F10192: entity F port map(lamdaA => P(10)(192),lamdaB => P(10)(193),lamdaOut => P(9)(192));
U_G10193: entity G port map(lamdaA => P(10)(192),lamdaB => P(10)(193),s => s(10)(96),lamdaOut => P(9)(193));
U_F10194: entity F port map(lamdaA => P(10)(194),lamdaB => P(10)(195),lamdaOut => P(9)(194));
U_G10195: entity G port map(lamdaA => P(10)(194),lamdaB => P(10)(195),s => s(10)(97),lamdaOut => P(9)(195));
U_F10196: entity F port map(lamdaA => P(10)(196),lamdaB => P(10)(197),lamdaOut => P(9)(196));
U_G10197: entity G port map(lamdaA => P(10)(196),lamdaB => P(10)(197),s => s(10)(98),lamdaOut => P(9)(197));
U_F10198: entity F port map(lamdaA => P(10)(198),lamdaB => P(10)(199),lamdaOut => P(9)(198));
U_G10199: entity G port map(lamdaA => P(10)(198),lamdaB => P(10)(199),s => s(10)(99),lamdaOut => P(9)(199));
U_F10200: entity F port map(lamdaA => P(10)(200),lamdaB => P(10)(201),lamdaOut => P(9)(200));
U_G10201: entity G port map(lamdaA => P(10)(200),lamdaB => P(10)(201),s => s(10)(100),lamdaOut => P(9)(201));
U_F10202: entity F port map(lamdaA => P(10)(202),lamdaB => P(10)(203),lamdaOut => P(9)(202));
U_G10203: entity G port map(lamdaA => P(10)(202),lamdaB => P(10)(203),s => s(10)(101),lamdaOut => P(9)(203));
U_F10204: entity F port map(lamdaA => P(10)(204),lamdaB => P(10)(205),lamdaOut => P(9)(204));
U_G10205: entity G port map(lamdaA => P(10)(204),lamdaB => P(10)(205),s => s(10)(102),lamdaOut => P(9)(205));
U_F10206: entity F port map(lamdaA => P(10)(206),lamdaB => P(10)(207),lamdaOut => P(9)(206));
U_G10207: entity G port map(lamdaA => P(10)(206),lamdaB => P(10)(207),s => s(10)(103),lamdaOut => P(9)(207));
U_F10208: entity F port map(lamdaA => P(10)(208),lamdaB => P(10)(209),lamdaOut => P(9)(208));
U_G10209: entity G port map(lamdaA => P(10)(208),lamdaB => P(10)(209),s => s(10)(104),lamdaOut => P(9)(209));
U_F10210: entity F port map(lamdaA => P(10)(210),lamdaB => P(10)(211),lamdaOut => P(9)(210));
U_G10211: entity G port map(lamdaA => P(10)(210),lamdaB => P(10)(211),s => s(10)(105),lamdaOut => P(9)(211));
U_F10212: entity F port map(lamdaA => P(10)(212),lamdaB => P(10)(213),lamdaOut => P(9)(212));
U_G10213: entity G port map(lamdaA => P(10)(212),lamdaB => P(10)(213),s => s(10)(106),lamdaOut => P(9)(213));
U_F10214: entity F port map(lamdaA => P(10)(214),lamdaB => P(10)(215),lamdaOut => P(9)(214));
U_G10215: entity G port map(lamdaA => P(10)(214),lamdaB => P(10)(215),s => s(10)(107),lamdaOut => P(9)(215));
U_F10216: entity F port map(lamdaA => P(10)(216),lamdaB => P(10)(217),lamdaOut => P(9)(216));
U_G10217: entity G port map(lamdaA => P(10)(216),lamdaB => P(10)(217),s => s(10)(108),lamdaOut => P(9)(217));
U_F10218: entity F port map(lamdaA => P(10)(218),lamdaB => P(10)(219),lamdaOut => P(9)(218));
U_G10219: entity G port map(lamdaA => P(10)(218),lamdaB => P(10)(219),s => s(10)(109),lamdaOut => P(9)(219));
U_F10220: entity F port map(lamdaA => P(10)(220),lamdaB => P(10)(221),lamdaOut => P(9)(220));
U_G10221: entity G port map(lamdaA => P(10)(220),lamdaB => P(10)(221),s => s(10)(110),lamdaOut => P(9)(221));
U_F10222: entity F port map(lamdaA => P(10)(222),lamdaB => P(10)(223),lamdaOut => P(9)(222));
U_G10223: entity G port map(lamdaA => P(10)(222),lamdaB => P(10)(223),s => s(10)(111),lamdaOut => P(9)(223));
U_F10224: entity F port map(lamdaA => P(10)(224),lamdaB => P(10)(225),lamdaOut => P(9)(224));
U_G10225: entity G port map(lamdaA => P(10)(224),lamdaB => P(10)(225),s => s(10)(112),lamdaOut => P(9)(225));
U_F10226: entity F port map(lamdaA => P(10)(226),lamdaB => P(10)(227),lamdaOut => P(9)(226));
U_G10227: entity G port map(lamdaA => P(10)(226),lamdaB => P(10)(227),s => s(10)(113),lamdaOut => P(9)(227));
U_F10228: entity F port map(lamdaA => P(10)(228),lamdaB => P(10)(229),lamdaOut => P(9)(228));
U_G10229: entity G port map(lamdaA => P(10)(228),lamdaB => P(10)(229),s => s(10)(114),lamdaOut => P(9)(229));
U_F10230: entity F port map(lamdaA => P(10)(230),lamdaB => P(10)(231),lamdaOut => P(9)(230));
U_G10231: entity G port map(lamdaA => P(10)(230),lamdaB => P(10)(231),s => s(10)(115),lamdaOut => P(9)(231));
U_F10232: entity F port map(lamdaA => P(10)(232),lamdaB => P(10)(233),lamdaOut => P(9)(232));
U_G10233: entity G port map(lamdaA => P(10)(232),lamdaB => P(10)(233),s => s(10)(116),lamdaOut => P(9)(233));
U_F10234: entity F port map(lamdaA => P(10)(234),lamdaB => P(10)(235),lamdaOut => P(9)(234));
U_G10235: entity G port map(lamdaA => P(10)(234),lamdaB => P(10)(235),s => s(10)(117),lamdaOut => P(9)(235));
U_F10236: entity F port map(lamdaA => P(10)(236),lamdaB => P(10)(237),lamdaOut => P(9)(236));
U_G10237: entity G port map(lamdaA => P(10)(236),lamdaB => P(10)(237),s => s(10)(118),lamdaOut => P(9)(237));
U_F10238: entity F port map(lamdaA => P(10)(238),lamdaB => P(10)(239),lamdaOut => P(9)(238));
U_G10239: entity G port map(lamdaA => P(10)(238),lamdaB => P(10)(239),s => s(10)(119),lamdaOut => P(9)(239));
U_F10240: entity F port map(lamdaA => P(10)(240),lamdaB => P(10)(241),lamdaOut => P(9)(240));
U_G10241: entity G port map(lamdaA => P(10)(240),lamdaB => P(10)(241),s => s(10)(120),lamdaOut => P(9)(241));
U_F10242: entity F port map(lamdaA => P(10)(242),lamdaB => P(10)(243),lamdaOut => P(9)(242));
U_G10243: entity G port map(lamdaA => P(10)(242),lamdaB => P(10)(243),s => s(10)(121),lamdaOut => P(9)(243));
U_F10244: entity F port map(lamdaA => P(10)(244),lamdaB => P(10)(245),lamdaOut => P(9)(244));
U_G10245: entity G port map(lamdaA => P(10)(244),lamdaB => P(10)(245),s => s(10)(122),lamdaOut => P(9)(245));
U_F10246: entity F port map(lamdaA => P(10)(246),lamdaB => P(10)(247),lamdaOut => P(9)(246));
U_G10247: entity G port map(lamdaA => P(10)(246),lamdaB => P(10)(247),s => s(10)(123),lamdaOut => P(9)(247));
U_F10248: entity F port map(lamdaA => P(10)(248),lamdaB => P(10)(249),lamdaOut => P(9)(248));
U_G10249: entity G port map(lamdaA => P(10)(248),lamdaB => P(10)(249),s => s(10)(124),lamdaOut => P(9)(249));
U_F10250: entity F port map(lamdaA => P(10)(250),lamdaB => P(10)(251),lamdaOut => P(9)(250));
U_G10251: entity G port map(lamdaA => P(10)(250),lamdaB => P(10)(251),s => s(10)(125),lamdaOut => P(9)(251));
U_F10252: entity F port map(lamdaA => P(10)(252),lamdaB => P(10)(253),lamdaOut => P(9)(252));
U_G10253: entity G port map(lamdaA => P(10)(252),lamdaB => P(10)(253),s => s(10)(126),lamdaOut => P(9)(253));
U_F10254: entity F port map(lamdaA => P(10)(254),lamdaB => P(10)(255),lamdaOut => P(9)(254));
U_G10255: entity G port map(lamdaA => P(10)(254),lamdaB => P(10)(255),s => s(10)(127),lamdaOut => P(9)(255));
U_F10256: entity F port map(lamdaA => P(10)(256),lamdaB => P(10)(257),lamdaOut => P(9)(256));
U_G10257: entity G port map(lamdaA => P(10)(256),lamdaB => P(10)(257),s => s(10)(128),lamdaOut => P(9)(257));
U_F10258: entity F port map(lamdaA => P(10)(258),lamdaB => P(10)(259),lamdaOut => P(9)(258));
U_G10259: entity G port map(lamdaA => P(10)(258),lamdaB => P(10)(259),s => s(10)(129),lamdaOut => P(9)(259));
U_F10260: entity F port map(lamdaA => P(10)(260),lamdaB => P(10)(261),lamdaOut => P(9)(260));
U_G10261: entity G port map(lamdaA => P(10)(260),lamdaB => P(10)(261),s => s(10)(130),lamdaOut => P(9)(261));
U_F10262: entity F port map(lamdaA => P(10)(262),lamdaB => P(10)(263),lamdaOut => P(9)(262));
U_G10263: entity G port map(lamdaA => P(10)(262),lamdaB => P(10)(263),s => s(10)(131),lamdaOut => P(9)(263));
U_F10264: entity F port map(lamdaA => P(10)(264),lamdaB => P(10)(265),lamdaOut => P(9)(264));
U_G10265: entity G port map(lamdaA => P(10)(264),lamdaB => P(10)(265),s => s(10)(132),lamdaOut => P(9)(265));
U_F10266: entity F port map(lamdaA => P(10)(266),lamdaB => P(10)(267),lamdaOut => P(9)(266));
U_G10267: entity G port map(lamdaA => P(10)(266),lamdaB => P(10)(267),s => s(10)(133),lamdaOut => P(9)(267));
U_F10268: entity F port map(lamdaA => P(10)(268),lamdaB => P(10)(269),lamdaOut => P(9)(268));
U_G10269: entity G port map(lamdaA => P(10)(268),lamdaB => P(10)(269),s => s(10)(134),lamdaOut => P(9)(269));
U_F10270: entity F port map(lamdaA => P(10)(270),lamdaB => P(10)(271),lamdaOut => P(9)(270));
U_G10271: entity G port map(lamdaA => P(10)(270),lamdaB => P(10)(271),s => s(10)(135),lamdaOut => P(9)(271));
U_F10272: entity F port map(lamdaA => P(10)(272),lamdaB => P(10)(273),lamdaOut => P(9)(272));
U_G10273: entity G port map(lamdaA => P(10)(272),lamdaB => P(10)(273),s => s(10)(136),lamdaOut => P(9)(273));
U_F10274: entity F port map(lamdaA => P(10)(274),lamdaB => P(10)(275),lamdaOut => P(9)(274));
U_G10275: entity G port map(lamdaA => P(10)(274),lamdaB => P(10)(275),s => s(10)(137),lamdaOut => P(9)(275));
U_F10276: entity F port map(lamdaA => P(10)(276),lamdaB => P(10)(277),lamdaOut => P(9)(276));
U_G10277: entity G port map(lamdaA => P(10)(276),lamdaB => P(10)(277),s => s(10)(138),lamdaOut => P(9)(277));
U_F10278: entity F port map(lamdaA => P(10)(278),lamdaB => P(10)(279),lamdaOut => P(9)(278));
U_G10279: entity G port map(lamdaA => P(10)(278),lamdaB => P(10)(279),s => s(10)(139),lamdaOut => P(9)(279));
U_F10280: entity F port map(lamdaA => P(10)(280),lamdaB => P(10)(281),lamdaOut => P(9)(280));
U_G10281: entity G port map(lamdaA => P(10)(280),lamdaB => P(10)(281),s => s(10)(140),lamdaOut => P(9)(281));
U_F10282: entity F port map(lamdaA => P(10)(282),lamdaB => P(10)(283),lamdaOut => P(9)(282));
U_G10283: entity G port map(lamdaA => P(10)(282),lamdaB => P(10)(283),s => s(10)(141),lamdaOut => P(9)(283));
U_F10284: entity F port map(lamdaA => P(10)(284),lamdaB => P(10)(285),lamdaOut => P(9)(284));
U_G10285: entity G port map(lamdaA => P(10)(284),lamdaB => P(10)(285),s => s(10)(142),lamdaOut => P(9)(285));
U_F10286: entity F port map(lamdaA => P(10)(286),lamdaB => P(10)(287),lamdaOut => P(9)(286));
U_G10287: entity G port map(lamdaA => P(10)(286),lamdaB => P(10)(287),s => s(10)(143),lamdaOut => P(9)(287));
U_F10288: entity F port map(lamdaA => P(10)(288),lamdaB => P(10)(289),lamdaOut => P(9)(288));
U_G10289: entity G port map(lamdaA => P(10)(288),lamdaB => P(10)(289),s => s(10)(144),lamdaOut => P(9)(289));
U_F10290: entity F port map(lamdaA => P(10)(290),lamdaB => P(10)(291),lamdaOut => P(9)(290));
U_G10291: entity G port map(lamdaA => P(10)(290),lamdaB => P(10)(291),s => s(10)(145),lamdaOut => P(9)(291));
U_F10292: entity F port map(lamdaA => P(10)(292),lamdaB => P(10)(293),lamdaOut => P(9)(292));
U_G10293: entity G port map(lamdaA => P(10)(292),lamdaB => P(10)(293),s => s(10)(146),lamdaOut => P(9)(293));
U_F10294: entity F port map(lamdaA => P(10)(294),lamdaB => P(10)(295),lamdaOut => P(9)(294));
U_G10295: entity G port map(lamdaA => P(10)(294),lamdaB => P(10)(295),s => s(10)(147),lamdaOut => P(9)(295));
U_F10296: entity F port map(lamdaA => P(10)(296),lamdaB => P(10)(297),lamdaOut => P(9)(296));
U_G10297: entity G port map(lamdaA => P(10)(296),lamdaB => P(10)(297),s => s(10)(148),lamdaOut => P(9)(297));
U_F10298: entity F port map(lamdaA => P(10)(298),lamdaB => P(10)(299),lamdaOut => P(9)(298));
U_G10299: entity G port map(lamdaA => P(10)(298),lamdaB => P(10)(299),s => s(10)(149),lamdaOut => P(9)(299));
U_F10300: entity F port map(lamdaA => P(10)(300),lamdaB => P(10)(301),lamdaOut => P(9)(300));
U_G10301: entity G port map(lamdaA => P(10)(300),lamdaB => P(10)(301),s => s(10)(150),lamdaOut => P(9)(301));
U_F10302: entity F port map(lamdaA => P(10)(302),lamdaB => P(10)(303),lamdaOut => P(9)(302));
U_G10303: entity G port map(lamdaA => P(10)(302),lamdaB => P(10)(303),s => s(10)(151),lamdaOut => P(9)(303));
U_F10304: entity F port map(lamdaA => P(10)(304),lamdaB => P(10)(305),lamdaOut => P(9)(304));
U_G10305: entity G port map(lamdaA => P(10)(304),lamdaB => P(10)(305),s => s(10)(152),lamdaOut => P(9)(305));
U_F10306: entity F port map(lamdaA => P(10)(306),lamdaB => P(10)(307),lamdaOut => P(9)(306));
U_G10307: entity G port map(lamdaA => P(10)(306),lamdaB => P(10)(307),s => s(10)(153),lamdaOut => P(9)(307));
U_F10308: entity F port map(lamdaA => P(10)(308),lamdaB => P(10)(309),lamdaOut => P(9)(308));
U_G10309: entity G port map(lamdaA => P(10)(308),lamdaB => P(10)(309),s => s(10)(154),lamdaOut => P(9)(309));
U_F10310: entity F port map(lamdaA => P(10)(310),lamdaB => P(10)(311),lamdaOut => P(9)(310));
U_G10311: entity G port map(lamdaA => P(10)(310),lamdaB => P(10)(311),s => s(10)(155),lamdaOut => P(9)(311));
U_F10312: entity F port map(lamdaA => P(10)(312),lamdaB => P(10)(313),lamdaOut => P(9)(312));
U_G10313: entity G port map(lamdaA => P(10)(312),lamdaB => P(10)(313),s => s(10)(156),lamdaOut => P(9)(313));
U_F10314: entity F port map(lamdaA => P(10)(314),lamdaB => P(10)(315),lamdaOut => P(9)(314));
U_G10315: entity G port map(lamdaA => P(10)(314),lamdaB => P(10)(315),s => s(10)(157),lamdaOut => P(9)(315));
U_F10316: entity F port map(lamdaA => P(10)(316),lamdaB => P(10)(317),lamdaOut => P(9)(316));
U_G10317: entity G port map(lamdaA => P(10)(316),lamdaB => P(10)(317),s => s(10)(158),lamdaOut => P(9)(317));
U_F10318: entity F port map(lamdaA => P(10)(318),lamdaB => P(10)(319),lamdaOut => P(9)(318));
U_G10319: entity G port map(lamdaA => P(10)(318),lamdaB => P(10)(319),s => s(10)(159),lamdaOut => P(9)(319));
U_F10320: entity F port map(lamdaA => P(10)(320),lamdaB => P(10)(321),lamdaOut => P(9)(320));
U_G10321: entity G port map(lamdaA => P(10)(320),lamdaB => P(10)(321),s => s(10)(160),lamdaOut => P(9)(321));
U_F10322: entity F port map(lamdaA => P(10)(322),lamdaB => P(10)(323),lamdaOut => P(9)(322));
U_G10323: entity G port map(lamdaA => P(10)(322),lamdaB => P(10)(323),s => s(10)(161),lamdaOut => P(9)(323));
U_F10324: entity F port map(lamdaA => P(10)(324),lamdaB => P(10)(325),lamdaOut => P(9)(324));
U_G10325: entity G port map(lamdaA => P(10)(324),lamdaB => P(10)(325),s => s(10)(162),lamdaOut => P(9)(325));
U_F10326: entity F port map(lamdaA => P(10)(326),lamdaB => P(10)(327),lamdaOut => P(9)(326));
U_G10327: entity G port map(lamdaA => P(10)(326),lamdaB => P(10)(327),s => s(10)(163),lamdaOut => P(9)(327));
U_F10328: entity F port map(lamdaA => P(10)(328),lamdaB => P(10)(329),lamdaOut => P(9)(328));
U_G10329: entity G port map(lamdaA => P(10)(328),lamdaB => P(10)(329),s => s(10)(164),lamdaOut => P(9)(329));
U_F10330: entity F port map(lamdaA => P(10)(330),lamdaB => P(10)(331),lamdaOut => P(9)(330));
U_G10331: entity G port map(lamdaA => P(10)(330),lamdaB => P(10)(331),s => s(10)(165),lamdaOut => P(9)(331));
U_F10332: entity F port map(lamdaA => P(10)(332),lamdaB => P(10)(333),lamdaOut => P(9)(332));
U_G10333: entity G port map(lamdaA => P(10)(332),lamdaB => P(10)(333),s => s(10)(166),lamdaOut => P(9)(333));
U_F10334: entity F port map(lamdaA => P(10)(334),lamdaB => P(10)(335),lamdaOut => P(9)(334));
U_G10335: entity G port map(lamdaA => P(10)(334),lamdaB => P(10)(335),s => s(10)(167),lamdaOut => P(9)(335));
U_F10336: entity F port map(lamdaA => P(10)(336),lamdaB => P(10)(337),lamdaOut => P(9)(336));
U_G10337: entity G port map(lamdaA => P(10)(336),lamdaB => P(10)(337),s => s(10)(168),lamdaOut => P(9)(337));
U_F10338: entity F port map(lamdaA => P(10)(338),lamdaB => P(10)(339),lamdaOut => P(9)(338));
U_G10339: entity G port map(lamdaA => P(10)(338),lamdaB => P(10)(339),s => s(10)(169),lamdaOut => P(9)(339));
U_F10340: entity F port map(lamdaA => P(10)(340),lamdaB => P(10)(341),lamdaOut => P(9)(340));
U_G10341: entity G port map(lamdaA => P(10)(340),lamdaB => P(10)(341),s => s(10)(170),lamdaOut => P(9)(341));
U_F10342: entity F port map(lamdaA => P(10)(342),lamdaB => P(10)(343),lamdaOut => P(9)(342));
U_G10343: entity G port map(lamdaA => P(10)(342),lamdaB => P(10)(343),s => s(10)(171),lamdaOut => P(9)(343));
U_F10344: entity F port map(lamdaA => P(10)(344),lamdaB => P(10)(345),lamdaOut => P(9)(344));
U_G10345: entity G port map(lamdaA => P(10)(344),lamdaB => P(10)(345),s => s(10)(172),lamdaOut => P(9)(345));
U_F10346: entity F port map(lamdaA => P(10)(346),lamdaB => P(10)(347),lamdaOut => P(9)(346));
U_G10347: entity G port map(lamdaA => P(10)(346),lamdaB => P(10)(347),s => s(10)(173),lamdaOut => P(9)(347));
U_F10348: entity F port map(lamdaA => P(10)(348),lamdaB => P(10)(349),lamdaOut => P(9)(348));
U_G10349: entity G port map(lamdaA => P(10)(348),lamdaB => P(10)(349),s => s(10)(174),lamdaOut => P(9)(349));
U_F10350: entity F port map(lamdaA => P(10)(350),lamdaB => P(10)(351),lamdaOut => P(9)(350));
U_G10351: entity G port map(lamdaA => P(10)(350),lamdaB => P(10)(351),s => s(10)(175),lamdaOut => P(9)(351));
U_F10352: entity F port map(lamdaA => P(10)(352),lamdaB => P(10)(353),lamdaOut => P(9)(352));
U_G10353: entity G port map(lamdaA => P(10)(352),lamdaB => P(10)(353),s => s(10)(176),lamdaOut => P(9)(353));
U_F10354: entity F port map(lamdaA => P(10)(354),lamdaB => P(10)(355),lamdaOut => P(9)(354));
U_G10355: entity G port map(lamdaA => P(10)(354),lamdaB => P(10)(355),s => s(10)(177),lamdaOut => P(9)(355));
U_F10356: entity F port map(lamdaA => P(10)(356),lamdaB => P(10)(357),lamdaOut => P(9)(356));
U_G10357: entity G port map(lamdaA => P(10)(356),lamdaB => P(10)(357),s => s(10)(178),lamdaOut => P(9)(357));
U_F10358: entity F port map(lamdaA => P(10)(358),lamdaB => P(10)(359),lamdaOut => P(9)(358));
U_G10359: entity G port map(lamdaA => P(10)(358),lamdaB => P(10)(359),s => s(10)(179),lamdaOut => P(9)(359));
U_F10360: entity F port map(lamdaA => P(10)(360),lamdaB => P(10)(361),lamdaOut => P(9)(360));
U_G10361: entity G port map(lamdaA => P(10)(360),lamdaB => P(10)(361),s => s(10)(180),lamdaOut => P(9)(361));
U_F10362: entity F port map(lamdaA => P(10)(362),lamdaB => P(10)(363),lamdaOut => P(9)(362));
U_G10363: entity G port map(lamdaA => P(10)(362),lamdaB => P(10)(363),s => s(10)(181),lamdaOut => P(9)(363));
U_F10364: entity F port map(lamdaA => P(10)(364),lamdaB => P(10)(365),lamdaOut => P(9)(364));
U_G10365: entity G port map(lamdaA => P(10)(364),lamdaB => P(10)(365),s => s(10)(182),lamdaOut => P(9)(365));
U_F10366: entity F port map(lamdaA => P(10)(366),lamdaB => P(10)(367),lamdaOut => P(9)(366));
U_G10367: entity G port map(lamdaA => P(10)(366),lamdaB => P(10)(367),s => s(10)(183),lamdaOut => P(9)(367));
U_F10368: entity F port map(lamdaA => P(10)(368),lamdaB => P(10)(369),lamdaOut => P(9)(368));
U_G10369: entity G port map(lamdaA => P(10)(368),lamdaB => P(10)(369),s => s(10)(184),lamdaOut => P(9)(369));
U_F10370: entity F port map(lamdaA => P(10)(370),lamdaB => P(10)(371),lamdaOut => P(9)(370));
U_G10371: entity G port map(lamdaA => P(10)(370),lamdaB => P(10)(371),s => s(10)(185),lamdaOut => P(9)(371));
U_F10372: entity F port map(lamdaA => P(10)(372),lamdaB => P(10)(373),lamdaOut => P(9)(372));
U_G10373: entity G port map(lamdaA => P(10)(372),lamdaB => P(10)(373),s => s(10)(186),lamdaOut => P(9)(373));
U_F10374: entity F port map(lamdaA => P(10)(374),lamdaB => P(10)(375),lamdaOut => P(9)(374));
U_G10375: entity G port map(lamdaA => P(10)(374),lamdaB => P(10)(375),s => s(10)(187),lamdaOut => P(9)(375));
U_F10376: entity F port map(lamdaA => P(10)(376),lamdaB => P(10)(377),lamdaOut => P(9)(376));
U_G10377: entity G port map(lamdaA => P(10)(376),lamdaB => P(10)(377),s => s(10)(188),lamdaOut => P(9)(377));
U_F10378: entity F port map(lamdaA => P(10)(378),lamdaB => P(10)(379),lamdaOut => P(9)(378));
U_G10379: entity G port map(lamdaA => P(10)(378),lamdaB => P(10)(379),s => s(10)(189),lamdaOut => P(9)(379));
U_F10380: entity F port map(lamdaA => P(10)(380),lamdaB => P(10)(381),lamdaOut => P(9)(380));
U_G10381: entity G port map(lamdaA => P(10)(380),lamdaB => P(10)(381),s => s(10)(190),lamdaOut => P(9)(381));
U_F10382: entity F port map(lamdaA => P(10)(382),lamdaB => P(10)(383),lamdaOut => P(9)(382));
U_G10383: entity G port map(lamdaA => P(10)(382),lamdaB => P(10)(383),s => s(10)(191),lamdaOut => P(9)(383));
U_F10384: entity F port map(lamdaA => P(10)(384),lamdaB => P(10)(385),lamdaOut => P(9)(384));
U_G10385: entity G port map(lamdaA => P(10)(384),lamdaB => P(10)(385),s => s(10)(192),lamdaOut => P(9)(385));
U_F10386: entity F port map(lamdaA => P(10)(386),lamdaB => P(10)(387),lamdaOut => P(9)(386));
U_G10387: entity G port map(lamdaA => P(10)(386),lamdaB => P(10)(387),s => s(10)(193),lamdaOut => P(9)(387));
U_F10388: entity F port map(lamdaA => P(10)(388),lamdaB => P(10)(389),lamdaOut => P(9)(388));
U_G10389: entity G port map(lamdaA => P(10)(388),lamdaB => P(10)(389),s => s(10)(194),lamdaOut => P(9)(389));
U_F10390: entity F port map(lamdaA => P(10)(390),lamdaB => P(10)(391),lamdaOut => P(9)(390));
U_G10391: entity G port map(lamdaA => P(10)(390),lamdaB => P(10)(391),s => s(10)(195),lamdaOut => P(9)(391));
U_F10392: entity F port map(lamdaA => P(10)(392),lamdaB => P(10)(393),lamdaOut => P(9)(392));
U_G10393: entity G port map(lamdaA => P(10)(392),lamdaB => P(10)(393),s => s(10)(196),lamdaOut => P(9)(393));
U_F10394: entity F port map(lamdaA => P(10)(394),lamdaB => P(10)(395),lamdaOut => P(9)(394));
U_G10395: entity G port map(lamdaA => P(10)(394),lamdaB => P(10)(395),s => s(10)(197),lamdaOut => P(9)(395));
U_F10396: entity F port map(lamdaA => P(10)(396),lamdaB => P(10)(397),lamdaOut => P(9)(396));
U_G10397: entity G port map(lamdaA => P(10)(396),lamdaB => P(10)(397),s => s(10)(198),lamdaOut => P(9)(397));
U_F10398: entity F port map(lamdaA => P(10)(398),lamdaB => P(10)(399),lamdaOut => P(9)(398));
U_G10399: entity G port map(lamdaA => P(10)(398),lamdaB => P(10)(399),s => s(10)(199),lamdaOut => P(9)(399));
U_F10400: entity F port map(lamdaA => P(10)(400),lamdaB => P(10)(401),lamdaOut => P(9)(400));
U_G10401: entity G port map(lamdaA => P(10)(400),lamdaB => P(10)(401),s => s(10)(200),lamdaOut => P(9)(401));
U_F10402: entity F port map(lamdaA => P(10)(402),lamdaB => P(10)(403),lamdaOut => P(9)(402));
U_G10403: entity G port map(lamdaA => P(10)(402),lamdaB => P(10)(403),s => s(10)(201),lamdaOut => P(9)(403));
U_F10404: entity F port map(lamdaA => P(10)(404),lamdaB => P(10)(405),lamdaOut => P(9)(404));
U_G10405: entity G port map(lamdaA => P(10)(404),lamdaB => P(10)(405),s => s(10)(202),lamdaOut => P(9)(405));
U_F10406: entity F port map(lamdaA => P(10)(406),lamdaB => P(10)(407),lamdaOut => P(9)(406));
U_G10407: entity G port map(lamdaA => P(10)(406),lamdaB => P(10)(407),s => s(10)(203),lamdaOut => P(9)(407));
U_F10408: entity F port map(lamdaA => P(10)(408),lamdaB => P(10)(409),lamdaOut => P(9)(408));
U_G10409: entity G port map(lamdaA => P(10)(408),lamdaB => P(10)(409),s => s(10)(204),lamdaOut => P(9)(409));
U_F10410: entity F port map(lamdaA => P(10)(410),lamdaB => P(10)(411),lamdaOut => P(9)(410));
U_G10411: entity G port map(lamdaA => P(10)(410),lamdaB => P(10)(411),s => s(10)(205),lamdaOut => P(9)(411));
U_F10412: entity F port map(lamdaA => P(10)(412),lamdaB => P(10)(413),lamdaOut => P(9)(412));
U_G10413: entity G port map(lamdaA => P(10)(412),lamdaB => P(10)(413),s => s(10)(206),lamdaOut => P(9)(413));
U_F10414: entity F port map(lamdaA => P(10)(414),lamdaB => P(10)(415),lamdaOut => P(9)(414));
U_G10415: entity G port map(lamdaA => P(10)(414),lamdaB => P(10)(415),s => s(10)(207),lamdaOut => P(9)(415));
U_F10416: entity F port map(lamdaA => P(10)(416),lamdaB => P(10)(417),lamdaOut => P(9)(416));
U_G10417: entity G port map(lamdaA => P(10)(416),lamdaB => P(10)(417),s => s(10)(208),lamdaOut => P(9)(417));
U_F10418: entity F port map(lamdaA => P(10)(418),lamdaB => P(10)(419),lamdaOut => P(9)(418));
U_G10419: entity G port map(lamdaA => P(10)(418),lamdaB => P(10)(419),s => s(10)(209),lamdaOut => P(9)(419));
U_F10420: entity F port map(lamdaA => P(10)(420),lamdaB => P(10)(421),lamdaOut => P(9)(420));
U_G10421: entity G port map(lamdaA => P(10)(420),lamdaB => P(10)(421),s => s(10)(210),lamdaOut => P(9)(421));
U_F10422: entity F port map(lamdaA => P(10)(422),lamdaB => P(10)(423),lamdaOut => P(9)(422));
U_G10423: entity G port map(lamdaA => P(10)(422),lamdaB => P(10)(423),s => s(10)(211),lamdaOut => P(9)(423));
U_F10424: entity F port map(lamdaA => P(10)(424),lamdaB => P(10)(425),lamdaOut => P(9)(424));
U_G10425: entity G port map(lamdaA => P(10)(424),lamdaB => P(10)(425),s => s(10)(212),lamdaOut => P(9)(425));
U_F10426: entity F port map(lamdaA => P(10)(426),lamdaB => P(10)(427),lamdaOut => P(9)(426));
U_G10427: entity G port map(lamdaA => P(10)(426),lamdaB => P(10)(427),s => s(10)(213),lamdaOut => P(9)(427));
U_F10428: entity F port map(lamdaA => P(10)(428),lamdaB => P(10)(429),lamdaOut => P(9)(428));
U_G10429: entity G port map(lamdaA => P(10)(428),lamdaB => P(10)(429),s => s(10)(214),lamdaOut => P(9)(429));
U_F10430: entity F port map(lamdaA => P(10)(430),lamdaB => P(10)(431),lamdaOut => P(9)(430));
U_G10431: entity G port map(lamdaA => P(10)(430),lamdaB => P(10)(431),s => s(10)(215),lamdaOut => P(9)(431));
U_F10432: entity F port map(lamdaA => P(10)(432),lamdaB => P(10)(433),lamdaOut => P(9)(432));
U_G10433: entity G port map(lamdaA => P(10)(432),lamdaB => P(10)(433),s => s(10)(216),lamdaOut => P(9)(433));
U_F10434: entity F port map(lamdaA => P(10)(434),lamdaB => P(10)(435),lamdaOut => P(9)(434));
U_G10435: entity G port map(lamdaA => P(10)(434),lamdaB => P(10)(435),s => s(10)(217),lamdaOut => P(9)(435));
U_F10436: entity F port map(lamdaA => P(10)(436),lamdaB => P(10)(437),lamdaOut => P(9)(436));
U_G10437: entity G port map(lamdaA => P(10)(436),lamdaB => P(10)(437),s => s(10)(218),lamdaOut => P(9)(437));
U_F10438: entity F port map(lamdaA => P(10)(438),lamdaB => P(10)(439),lamdaOut => P(9)(438));
U_G10439: entity G port map(lamdaA => P(10)(438),lamdaB => P(10)(439),s => s(10)(219),lamdaOut => P(9)(439));
U_F10440: entity F port map(lamdaA => P(10)(440),lamdaB => P(10)(441),lamdaOut => P(9)(440));
U_G10441: entity G port map(lamdaA => P(10)(440),lamdaB => P(10)(441),s => s(10)(220),lamdaOut => P(9)(441));
U_F10442: entity F port map(lamdaA => P(10)(442),lamdaB => P(10)(443),lamdaOut => P(9)(442));
U_G10443: entity G port map(lamdaA => P(10)(442),lamdaB => P(10)(443),s => s(10)(221),lamdaOut => P(9)(443));
U_F10444: entity F port map(lamdaA => P(10)(444),lamdaB => P(10)(445),lamdaOut => P(9)(444));
U_G10445: entity G port map(lamdaA => P(10)(444),lamdaB => P(10)(445),s => s(10)(222),lamdaOut => P(9)(445));
U_F10446: entity F port map(lamdaA => P(10)(446),lamdaB => P(10)(447),lamdaOut => P(9)(446));
U_G10447: entity G port map(lamdaA => P(10)(446),lamdaB => P(10)(447),s => s(10)(223),lamdaOut => P(9)(447));
U_F10448: entity F port map(lamdaA => P(10)(448),lamdaB => P(10)(449),lamdaOut => P(9)(448));
U_G10449: entity G port map(lamdaA => P(10)(448),lamdaB => P(10)(449),s => s(10)(224),lamdaOut => P(9)(449));
U_F10450: entity F port map(lamdaA => P(10)(450),lamdaB => P(10)(451),lamdaOut => P(9)(450));
U_G10451: entity G port map(lamdaA => P(10)(450),lamdaB => P(10)(451),s => s(10)(225),lamdaOut => P(9)(451));
U_F10452: entity F port map(lamdaA => P(10)(452),lamdaB => P(10)(453),lamdaOut => P(9)(452));
U_G10453: entity G port map(lamdaA => P(10)(452),lamdaB => P(10)(453),s => s(10)(226),lamdaOut => P(9)(453));
U_F10454: entity F port map(lamdaA => P(10)(454),lamdaB => P(10)(455),lamdaOut => P(9)(454));
U_G10455: entity G port map(lamdaA => P(10)(454),lamdaB => P(10)(455),s => s(10)(227),lamdaOut => P(9)(455));
U_F10456: entity F port map(lamdaA => P(10)(456),lamdaB => P(10)(457),lamdaOut => P(9)(456));
U_G10457: entity G port map(lamdaA => P(10)(456),lamdaB => P(10)(457),s => s(10)(228),lamdaOut => P(9)(457));
U_F10458: entity F port map(lamdaA => P(10)(458),lamdaB => P(10)(459),lamdaOut => P(9)(458));
U_G10459: entity G port map(lamdaA => P(10)(458),lamdaB => P(10)(459),s => s(10)(229),lamdaOut => P(9)(459));
U_F10460: entity F port map(lamdaA => P(10)(460),lamdaB => P(10)(461),lamdaOut => P(9)(460));
U_G10461: entity G port map(lamdaA => P(10)(460),lamdaB => P(10)(461),s => s(10)(230),lamdaOut => P(9)(461));
U_F10462: entity F port map(lamdaA => P(10)(462),lamdaB => P(10)(463),lamdaOut => P(9)(462));
U_G10463: entity G port map(lamdaA => P(10)(462),lamdaB => P(10)(463),s => s(10)(231),lamdaOut => P(9)(463));
U_F10464: entity F port map(lamdaA => P(10)(464),lamdaB => P(10)(465),lamdaOut => P(9)(464));
U_G10465: entity G port map(lamdaA => P(10)(464),lamdaB => P(10)(465),s => s(10)(232),lamdaOut => P(9)(465));
U_F10466: entity F port map(lamdaA => P(10)(466),lamdaB => P(10)(467),lamdaOut => P(9)(466));
U_G10467: entity G port map(lamdaA => P(10)(466),lamdaB => P(10)(467),s => s(10)(233),lamdaOut => P(9)(467));
U_F10468: entity F port map(lamdaA => P(10)(468),lamdaB => P(10)(469),lamdaOut => P(9)(468));
U_G10469: entity G port map(lamdaA => P(10)(468),lamdaB => P(10)(469),s => s(10)(234),lamdaOut => P(9)(469));
U_F10470: entity F port map(lamdaA => P(10)(470),lamdaB => P(10)(471),lamdaOut => P(9)(470));
U_G10471: entity G port map(lamdaA => P(10)(470),lamdaB => P(10)(471),s => s(10)(235),lamdaOut => P(9)(471));
U_F10472: entity F port map(lamdaA => P(10)(472),lamdaB => P(10)(473),lamdaOut => P(9)(472));
U_G10473: entity G port map(lamdaA => P(10)(472),lamdaB => P(10)(473),s => s(10)(236),lamdaOut => P(9)(473));
U_F10474: entity F port map(lamdaA => P(10)(474),lamdaB => P(10)(475),lamdaOut => P(9)(474));
U_G10475: entity G port map(lamdaA => P(10)(474),lamdaB => P(10)(475),s => s(10)(237),lamdaOut => P(9)(475));
U_F10476: entity F port map(lamdaA => P(10)(476),lamdaB => P(10)(477),lamdaOut => P(9)(476));
U_G10477: entity G port map(lamdaA => P(10)(476),lamdaB => P(10)(477),s => s(10)(238),lamdaOut => P(9)(477));
U_F10478: entity F port map(lamdaA => P(10)(478),lamdaB => P(10)(479),lamdaOut => P(9)(478));
U_G10479: entity G port map(lamdaA => P(10)(478),lamdaB => P(10)(479),s => s(10)(239),lamdaOut => P(9)(479));
U_F10480: entity F port map(lamdaA => P(10)(480),lamdaB => P(10)(481),lamdaOut => P(9)(480));
U_G10481: entity G port map(lamdaA => P(10)(480),lamdaB => P(10)(481),s => s(10)(240),lamdaOut => P(9)(481));
U_F10482: entity F port map(lamdaA => P(10)(482),lamdaB => P(10)(483),lamdaOut => P(9)(482));
U_G10483: entity G port map(lamdaA => P(10)(482),lamdaB => P(10)(483),s => s(10)(241),lamdaOut => P(9)(483));
U_F10484: entity F port map(lamdaA => P(10)(484),lamdaB => P(10)(485),lamdaOut => P(9)(484));
U_G10485: entity G port map(lamdaA => P(10)(484),lamdaB => P(10)(485),s => s(10)(242),lamdaOut => P(9)(485));
U_F10486: entity F port map(lamdaA => P(10)(486),lamdaB => P(10)(487),lamdaOut => P(9)(486));
U_G10487: entity G port map(lamdaA => P(10)(486),lamdaB => P(10)(487),s => s(10)(243),lamdaOut => P(9)(487));
U_F10488: entity F port map(lamdaA => P(10)(488),lamdaB => P(10)(489),lamdaOut => P(9)(488));
U_G10489: entity G port map(lamdaA => P(10)(488),lamdaB => P(10)(489),s => s(10)(244),lamdaOut => P(9)(489));
U_F10490: entity F port map(lamdaA => P(10)(490),lamdaB => P(10)(491),lamdaOut => P(9)(490));
U_G10491: entity G port map(lamdaA => P(10)(490),lamdaB => P(10)(491),s => s(10)(245),lamdaOut => P(9)(491));
U_F10492: entity F port map(lamdaA => P(10)(492),lamdaB => P(10)(493),lamdaOut => P(9)(492));
U_G10493: entity G port map(lamdaA => P(10)(492),lamdaB => P(10)(493),s => s(10)(246),lamdaOut => P(9)(493));
U_F10494: entity F port map(lamdaA => P(10)(494),lamdaB => P(10)(495),lamdaOut => P(9)(494));
U_G10495: entity G port map(lamdaA => P(10)(494),lamdaB => P(10)(495),s => s(10)(247),lamdaOut => P(9)(495));
U_F10496: entity F port map(lamdaA => P(10)(496),lamdaB => P(10)(497),lamdaOut => P(9)(496));
U_G10497: entity G port map(lamdaA => P(10)(496),lamdaB => P(10)(497),s => s(10)(248),lamdaOut => P(9)(497));
U_F10498: entity F port map(lamdaA => P(10)(498),lamdaB => P(10)(499),lamdaOut => P(9)(498));
U_G10499: entity G port map(lamdaA => P(10)(498),lamdaB => P(10)(499),s => s(10)(249),lamdaOut => P(9)(499));
U_F10500: entity F port map(lamdaA => P(10)(500),lamdaB => P(10)(501),lamdaOut => P(9)(500));
U_G10501: entity G port map(lamdaA => P(10)(500),lamdaB => P(10)(501),s => s(10)(250),lamdaOut => P(9)(501));
U_F10502: entity F port map(lamdaA => P(10)(502),lamdaB => P(10)(503),lamdaOut => P(9)(502));
U_G10503: entity G port map(lamdaA => P(10)(502),lamdaB => P(10)(503),s => s(10)(251),lamdaOut => P(9)(503));
U_F10504: entity F port map(lamdaA => P(10)(504),lamdaB => P(10)(505),lamdaOut => P(9)(504));
U_G10505: entity G port map(lamdaA => P(10)(504),lamdaB => P(10)(505),s => s(10)(252),lamdaOut => P(9)(505));
U_F10506: entity F port map(lamdaA => P(10)(506),lamdaB => P(10)(507),lamdaOut => P(9)(506));
U_G10507: entity G port map(lamdaA => P(10)(506),lamdaB => P(10)(507),s => s(10)(253),lamdaOut => P(9)(507));
U_F10508: entity F port map(lamdaA => P(10)(508),lamdaB => P(10)(509),lamdaOut => P(9)(508));
U_G10509: entity G port map(lamdaA => P(10)(508),lamdaB => P(10)(509),s => s(10)(254),lamdaOut => P(9)(509));
U_F10510: entity F port map(lamdaA => P(10)(510),lamdaB => P(10)(511),lamdaOut => P(9)(510));
U_G10511: entity G port map(lamdaA => P(10)(510),lamdaB => P(10)(511),s => s(10)(255),lamdaOut => P(9)(511));
U_F10512: entity F port map(lamdaA => P(10)(512),lamdaB => P(10)(513),lamdaOut => P(9)(512));
U_G10513: entity G port map(lamdaA => P(10)(512),lamdaB => P(10)(513),s => s(10)(256),lamdaOut => P(9)(513));
U_F10514: entity F port map(lamdaA => P(10)(514),lamdaB => P(10)(515),lamdaOut => P(9)(514));
U_G10515: entity G port map(lamdaA => P(10)(514),lamdaB => P(10)(515),s => s(10)(257),lamdaOut => P(9)(515));
U_F10516: entity F port map(lamdaA => P(10)(516),lamdaB => P(10)(517),lamdaOut => P(9)(516));
U_G10517: entity G port map(lamdaA => P(10)(516),lamdaB => P(10)(517),s => s(10)(258),lamdaOut => P(9)(517));
U_F10518: entity F port map(lamdaA => P(10)(518),lamdaB => P(10)(519),lamdaOut => P(9)(518));
U_G10519: entity G port map(lamdaA => P(10)(518),lamdaB => P(10)(519),s => s(10)(259),lamdaOut => P(9)(519));
U_F10520: entity F port map(lamdaA => P(10)(520),lamdaB => P(10)(521),lamdaOut => P(9)(520));
U_G10521: entity G port map(lamdaA => P(10)(520),lamdaB => P(10)(521),s => s(10)(260),lamdaOut => P(9)(521));
U_F10522: entity F port map(lamdaA => P(10)(522),lamdaB => P(10)(523),lamdaOut => P(9)(522));
U_G10523: entity G port map(lamdaA => P(10)(522),lamdaB => P(10)(523),s => s(10)(261),lamdaOut => P(9)(523));
U_F10524: entity F port map(lamdaA => P(10)(524),lamdaB => P(10)(525),lamdaOut => P(9)(524));
U_G10525: entity G port map(lamdaA => P(10)(524),lamdaB => P(10)(525),s => s(10)(262),lamdaOut => P(9)(525));
U_F10526: entity F port map(lamdaA => P(10)(526),lamdaB => P(10)(527),lamdaOut => P(9)(526));
U_G10527: entity G port map(lamdaA => P(10)(526),lamdaB => P(10)(527),s => s(10)(263),lamdaOut => P(9)(527));
U_F10528: entity F port map(lamdaA => P(10)(528),lamdaB => P(10)(529),lamdaOut => P(9)(528));
U_G10529: entity G port map(lamdaA => P(10)(528),lamdaB => P(10)(529),s => s(10)(264),lamdaOut => P(9)(529));
U_F10530: entity F port map(lamdaA => P(10)(530),lamdaB => P(10)(531),lamdaOut => P(9)(530));
U_G10531: entity G port map(lamdaA => P(10)(530),lamdaB => P(10)(531),s => s(10)(265),lamdaOut => P(9)(531));
U_F10532: entity F port map(lamdaA => P(10)(532),lamdaB => P(10)(533),lamdaOut => P(9)(532));
U_G10533: entity G port map(lamdaA => P(10)(532),lamdaB => P(10)(533),s => s(10)(266),lamdaOut => P(9)(533));
U_F10534: entity F port map(lamdaA => P(10)(534),lamdaB => P(10)(535),lamdaOut => P(9)(534));
U_G10535: entity G port map(lamdaA => P(10)(534),lamdaB => P(10)(535),s => s(10)(267),lamdaOut => P(9)(535));
U_F10536: entity F port map(lamdaA => P(10)(536),lamdaB => P(10)(537),lamdaOut => P(9)(536));
U_G10537: entity G port map(lamdaA => P(10)(536),lamdaB => P(10)(537),s => s(10)(268),lamdaOut => P(9)(537));
U_F10538: entity F port map(lamdaA => P(10)(538),lamdaB => P(10)(539),lamdaOut => P(9)(538));
U_G10539: entity G port map(lamdaA => P(10)(538),lamdaB => P(10)(539),s => s(10)(269),lamdaOut => P(9)(539));
U_F10540: entity F port map(lamdaA => P(10)(540),lamdaB => P(10)(541),lamdaOut => P(9)(540));
U_G10541: entity G port map(lamdaA => P(10)(540),lamdaB => P(10)(541),s => s(10)(270),lamdaOut => P(9)(541));
U_F10542: entity F port map(lamdaA => P(10)(542),lamdaB => P(10)(543),lamdaOut => P(9)(542));
U_G10543: entity G port map(lamdaA => P(10)(542),lamdaB => P(10)(543),s => s(10)(271),lamdaOut => P(9)(543));
U_F10544: entity F port map(lamdaA => P(10)(544),lamdaB => P(10)(545),lamdaOut => P(9)(544));
U_G10545: entity G port map(lamdaA => P(10)(544),lamdaB => P(10)(545),s => s(10)(272),lamdaOut => P(9)(545));
U_F10546: entity F port map(lamdaA => P(10)(546),lamdaB => P(10)(547),lamdaOut => P(9)(546));
U_G10547: entity G port map(lamdaA => P(10)(546),lamdaB => P(10)(547),s => s(10)(273),lamdaOut => P(9)(547));
U_F10548: entity F port map(lamdaA => P(10)(548),lamdaB => P(10)(549),lamdaOut => P(9)(548));
U_G10549: entity G port map(lamdaA => P(10)(548),lamdaB => P(10)(549),s => s(10)(274),lamdaOut => P(9)(549));
U_F10550: entity F port map(lamdaA => P(10)(550),lamdaB => P(10)(551),lamdaOut => P(9)(550));
U_G10551: entity G port map(lamdaA => P(10)(550),lamdaB => P(10)(551),s => s(10)(275),lamdaOut => P(9)(551));
U_F10552: entity F port map(lamdaA => P(10)(552),lamdaB => P(10)(553),lamdaOut => P(9)(552));
U_G10553: entity G port map(lamdaA => P(10)(552),lamdaB => P(10)(553),s => s(10)(276),lamdaOut => P(9)(553));
U_F10554: entity F port map(lamdaA => P(10)(554),lamdaB => P(10)(555),lamdaOut => P(9)(554));
U_G10555: entity G port map(lamdaA => P(10)(554),lamdaB => P(10)(555),s => s(10)(277),lamdaOut => P(9)(555));
U_F10556: entity F port map(lamdaA => P(10)(556),lamdaB => P(10)(557),lamdaOut => P(9)(556));
U_G10557: entity G port map(lamdaA => P(10)(556),lamdaB => P(10)(557),s => s(10)(278),lamdaOut => P(9)(557));
U_F10558: entity F port map(lamdaA => P(10)(558),lamdaB => P(10)(559),lamdaOut => P(9)(558));
U_G10559: entity G port map(lamdaA => P(10)(558),lamdaB => P(10)(559),s => s(10)(279),lamdaOut => P(9)(559));
U_F10560: entity F port map(lamdaA => P(10)(560),lamdaB => P(10)(561),lamdaOut => P(9)(560));
U_G10561: entity G port map(lamdaA => P(10)(560),lamdaB => P(10)(561),s => s(10)(280),lamdaOut => P(9)(561));
U_F10562: entity F port map(lamdaA => P(10)(562),lamdaB => P(10)(563),lamdaOut => P(9)(562));
U_G10563: entity G port map(lamdaA => P(10)(562),lamdaB => P(10)(563),s => s(10)(281),lamdaOut => P(9)(563));
U_F10564: entity F port map(lamdaA => P(10)(564),lamdaB => P(10)(565),lamdaOut => P(9)(564));
U_G10565: entity G port map(lamdaA => P(10)(564),lamdaB => P(10)(565),s => s(10)(282),lamdaOut => P(9)(565));
U_F10566: entity F port map(lamdaA => P(10)(566),lamdaB => P(10)(567),lamdaOut => P(9)(566));
U_G10567: entity G port map(lamdaA => P(10)(566),lamdaB => P(10)(567),s => s(10)(283),lamdaOut => P(9)(567));
U_F10568: entity F port map(lamdaA => P(10)(568),lamdaB => P(10)(569),lamdaOut => P(9)(568));
U_G10569: entity G port map(lamdaA => P(10)(568),lamdaB => P(10)(569),s => s(10)(284),lamdaOut => P(9)(569));
U_F10570: entity F port map(lamdaA => P(10)(570),lamdaB => P(10)(571),lamdaOut => P(9)(570));
U_G10571: entity G port map(lamdaA => P(10)(570),lamdaB => P(10)(571),s => s(10)(285),lamdaOut => P(9)(571));
U_F10572: entity F port map(lamdaA => P(10)(572),lamdaB => P(10)(573),lamdaOut => P(9)(572));
U_G10573: entity G port map(lamdaA => P(10)(572),lamdaB => P(10)(573),s => s(10)(286),lamdaOut => P(9)(573));
U_F10574: entity F port map(lamdaA => P(10)(574),lamdaB => P(10)(575),lamdaOut => P(9)(574));
U_G10575: entity G port map(lamdaA => P(10)(574),lamdaB => P(10)(575),s => s(10)(287),lamdaOut => P(9)(575));
U_F10576: entity F port map(lamdaA => P(10)(576),lamdaB => P(10)(577),lamdaOut => P(9)(576));
U_G10577: entity G port map(lamdaA => P(10)(576),lamdaB => P(10)(577),s => s(10)(288),lamdaOut => P(9)(577));
U_F10578: entity F port map(lamdaA => P(10)(578),lamdaB => P(10)(579),lamdaOut => P(9)(578));
U_G10579: entity G port map(lamdaA => P(10)(578),lamdaB => P(10)(579),s => s(10)(289),lamdaOut => P(9)(579));
U_F10580: entity F port map(lamdaA => P(10)(580),lamdaB => P(10)(581),lamdaOut => P(9)(580));
U_G10581: entity G port map(lamdaA => P(10)(580),lamdaB => P(10)(581),s => s(10)(290),lamdaOut => P(9)(581));
U_F10582: entity F port map(lamdaA => P(10)(582),lamdaB => P(10)(583),lamdaOut => P(9)(582));
U_G10583: entity G port map(lamdaA => P(10)(582),lamdaB => P(10)(583),s => s(10)(291),lamdaOut => P(9)(583));
U_F10584: entity F port map(lamdaA => P(10)(584),lamdaB => P(10)(585),lamdaOut => P(9)(584));
U_G10585: entity G port map(lamdaA => P(10)(584),lamdaB => P(10)(585),s => s(10)(292),lamdaOut => P(9)(585));
U_F10586: entity F port map(lamdaA => P(10)(586),lamdaB => P(10)(587),lamdaOut => P(9)(586));
U_G10587: entity G port map(lamdaA => P(10)(586),lamdaB => P(10)(587),s => s(10)(293),lamdaOut => P(9)(587));
U_F10588: entity F port map(lamdaA => P(10)(588),lamdaB => P(10)(589),lamdaOut => P(9)(588));
U_G10589: entity G port map(lamdaA => P(10)(588),lamdaB => P(10)(589),s => s(10)(294),lamdaOut => P(9)(589));
U_F10590: entity F port map(lamdaA => P(10)(590),lamdaB => P(10)(591),lamdaOut => P(9)(590));
U_G10591: entity G port map(lamdaA => P(10)(590),lamdaB => P(10)(591),s => s(10)(295),lamdaOut => P(9)(591));
U_F10592: entity F port map(lamdaA => P(10)(592),lamdaB => P(10)(593),lamdaOut => P(9)(592));
U_G10593: entity G port map(lamdaA => P(10)(592),lamdaB => P(10)(593),s => s(10)(296),lamdaOut => P(9)(593));
U_F10594: entity F port map(lamdaA => P(10)(594),lamdaB => P(10)(595),lamdaOut => P(9)(594));
U_G10595: entity G port map(lamdaA => P(10)(594),lamdaB => P(10)(595),s => s(10)(297),lamdaOut => P(9)(595));
U_F10596: entity F port map(lamdaA => P(10)(596),lamdaB => P(10)(597),lamdaOut => P(9)(596));
U_G10597: entity G port map(lamdaA => P(10)(596),lamdaB => P(10)(597),s => s(10)(298),lamdaOut => P(9)(597));
U_F10598: entity F port map(lamdaA => P(10)(598),lamdaB => P(10)(599),lamdaOut => P(9)(598));
U_G10599: entity G port map(lamdaA => P(10)(598),lamdaB => P(10)(599),s => s(10)(299),lamdaOut => P(9)(599));
U_F10600: entity F port map(lamdaA => P(10)(600),lamdaB => P(10)(601),lamdaOut => P(9)(600));
U_G10601: entity G port map(lamdaA => P(10)(600),lamdaB => P(10)(601),s => s(10)(300),lamdaOut => P(9)(601));
U_F10602: entity F port map(lamdaA => P(10)(602),lamdaB => P(10)(603),lamdaOut => P(9)(602));
U_G10603: entity G port map(lamdaA => P(10)(602),lamdaB => P(10)(603),s => s(10)(301),lamdaOut => P(9)(603));
U_F10604: entity F port map(lamdaA => P(10)(604),lamdaB => P(10)(605),lamdaOut => P(9)(604));
U_G10605: entity G port map(lamdaA => P(10)(604),lamdaB => P(10)(605),s => s(10)(302),lamdaOut => P(9)(605));
U_F10606: entity F port map(lamdaA => P(10)(606),lamdaB => P(10)(607),lamdaOut => P(9)(606));
U_G10607: entity G port map(lamdaA => P(10)(606),lamdaB => P(10)(607),s => s(10)(303),lamdaOut => P(9)(607));
U_F10608: entity F port map(lamdaA => P(10)(608),lamdaB => P(10)(609),lamdaOut => P(9)(608));
U_G10609: entity G port map(lamdaA => P(10)(608),lamdaB => P(10)(609),s => s(10)(304),lamdaOut => P(9)(609));
U_F10610: entity F port map(lamdaA => P(10)(610),lamdaB => P(10)(611),lamdaOut => P(9)(610));
U_G10611: entity G port map(lamdaA => P(10)(610),lamdaB => P(10)(611),s => s(10)(305),lamdaOut => P(9)(611));
U_F10612: entity F port map(lamdaA => P(10)(612),lamdaB => P(10)(613),lamdaOut => P(9)(612));
U_G10613: entity G port map(lamdaA => P(10)(612),lamdaB => P(10)(613),s => s(10)(306),lamdaOut => P(9)(613));
U_F10614: entity F port map(lamdaA => P(10)(614),lamdaB => P(10)(615),lamdaOut => P(9)(614));
U_G10615: entity G port map(lamdaA => P(10)(614),lamdaB => P(10)(615),s => s(10)(307),lamdaOut => P(9)(615));
U_F10616: entity F port map(lamdaA => P(10)(616),lamdaB => P(10)(617),lamdaOut => P(9)(616));
U_G10617: entity G port map(lamdaA => P(10)(616),lamdaB => P(10)(617),s => s(10)(308),lamdaOut => P(9)(617));
U_F10618: entity F port map(lamdaA => P(10)(618),lamdaB => P(10)(619),lamdaOut => P(9)(618));
U_G10619: entity G port map(lamdaA => P(10)(618),lamdaB => P(10)(619),s => s(10)(309),lamdaOut => P(9)(619));
U_F10620: entity F port map(lamdaA => P(10)(620),lamdaB => P(10)(621),lamdaOut => P(9)(620));
U_G10621: entity G port map(lamdaA => P(10)(620),lamdaB => P(10)(621),s => s(10)(310),lamdaOut => P(9)(621));
U_F10622: entity F port map(lamdaA => P(10)(622),lamdaB => P(10)(623),lamdaOut => P(9)(622));
U_G10623: entity G port map(lamdaA => P(10)(622),lamdaB => P(10)(623),s => s(10)(311),lamdaOut => P(9)(623));
U_F10624: entity F port map(lamdaA => P(10)(624),lamdaB => P(10)(625),lamdaOut => P(9)(624));
U_G10625: entity G port map(lamdaA => P(10)(624),lamdaB => P(10)(625),s => s(10)(312),lamdaOut => P(9)(625));
U_F10626: entity F port map(lamdaA => P(10)(626),lamdaB => P(10)(627),lamdaOut => P(9)(626));
U_G10627: entity G port map(lamdaA => P(10)(626),lamdaB => P(10)(627),s => s(10)(313),lamdaOut => P(9)(627));
U_F10628: entity F port map(lamdaA => P(10)(628),lamdaB => P(10)(629),lamdaOut => P(9)(628));
U_G10629: entity G port map(lamdaA => P(10)(628),lamdaB => P(10)(629),s => s(10)(314),lamdaOut => P(9)(629));
U_F10630: entity F port map(lamdaA => P(10)(630),lamdaB => P(10)(631),lamdaOut => P(9)(630));
U_G10631: entity G port map(lamdaA => P(10)(630),lamdaB => P(10)(631),s => s(10)(315),lamdaOut => P(9)(631));
U_F10632: entity F port map(lamdaA => P(10)(632),lamdaB => P(10)(633),lamdaOut => P(9)(632));
U_G10633: entity G port map(lamdaA => P(10)(632),lamdaB => P(10)(633),s => s(10)(316),lamdaOut => P(9)(633));
U_F10634: entity F port map(lamdaA => P(10)(634),lamdaB => P(10)(635),lamdaOut => P(9)(634));
U_G10635: entity G port map(lamdaA => P(10)(634),lamdaB => P(10)(635),s => s(10)(317),lamdaOut => P(9)(635));
U_F10636: entity F port map(lamdaA => P(10)(636),lamdaB => P(10)(637),lamdaOut => P(9)(636));
U_G10637: entity G port map(lamdaA => P(10)(636),lamdaB => P(10)(637),s => s(10)(318),lamdaOut => P(9)(637));
U_F10638: entity F port map(lamdaA => P(10)(638),lamdaB => P(10)(639),lamdaOut => P(9)(638));
U_G10639: entity G port map(lamdaA => P(10)(638),lamdaB => P(10)(639),s => s(10)(319),lamdaOut => P(9)(639));
U_F10640: entity F port map(lamdaA => P(10)(640),lamdaB => P(10)(641),lamdaOut => P(9)(640));
U_G10641: entity G port map(lamdaA => P(10)(640),lamdaB => P(10)(641),s => s(10)(320),lamdaOut => P(9)(641));
U_F10642: entity F port map(lamdaA => P(10)(642),lamdaB => P(10)(643),lamdaOut => P(9)(642));
U_G10643: entity G port map(lamdaA => P(10)(642),lamdaB => P(10)(643),s => s(10)(321),lamdaOut => P(9)(643));
U_F10644: entity F port map(lamdaA => P(10)(644),lamdaB => P(10)(645),lamdaOut => P(9)(644));
U_G10645: entity G port map(lamdaA => P(10)(644),lamdaB => P(10)(645),s => s(10)(322),lamdaOut => P(9)(645));
U_F10646: entity F port map(lamdaA => P(10)(646),lamdaB => P(10)(647),lamdaOut => P(9)(646));
U_G10647: entity G port map(lamdaA => P(10)(646),lamdaB => P(10)(647),s => s(10)(323),lamdaOut => P(9)(647));
U_F10648: entity F port map(lamdaA => P(10)(648),lamdaB => P(10)(649),lamdaOut => P(9)(648));
U_G10649: entity G port map(lamdaA => P(10)(648),lamdaB => P(10)(649),s => s(10)(324),lamdaOut => P(9)(649));
U_F10650: entity F port map(lamdaA => P(10)(650),lamdaB => P(10)(651),lamdaOut => P(9)(650));
U_G10651: entity G port map(lamdaA => P(10)(650),lamdaB => P(10)(651),s => s(10)(325),lamdaOut => P(9)(651));
U_F10652: entity F port map(lamdaA => P(10)(652),lamdaB => P(10)(653),lamdaOut => P(9)(652));
U_G10653: entity G port map(lamdaA => P(10)(652),lamdaB => P(10)(653),s => s(10)(326),lamdaOut => P(9)(653));
U_F10654: entity F port map(lamdaA => P(10)(654),lamdaB => P(10)(655),lamdaOut => P(9)(654));
U_G10655: entity G port map(lamdaA => P(10)(654),lamdaB => P(10)(655),s => s(10)(327),lamdaOut => P(9)(655));
U_F10656: entity F port map(lamdaA => P(10)(656),lamdaB => P(10)(657),lamdaOut => P(9)(656));
U_G10657: entity G port map(lamdaA => P(10)(656),lamdaB => P(10)(657),s => s(10)(328),lamdaOut => P(9)(657));
U_F10658: entity F port map(lamdaA => P(10)(658),lamdaB => P(10)(659),lamdaOut => P(9)(658));
U_G10659: entity G port map(lamdaA => P(10)(658),lamdaB => P(10)(659),s => s(10)(329),lamdaOut => P(9)(659));
U_F10660: entity F port map(lamdaA => P(10)(660),lamdaB => P(10)(661),lamdaOut => P(9)(660));
U_G10661: entity G port map(lamdaA => P(10)(660),lamdaB => P(10)(661),s => s(10)(330),lamdaOut => P(9)(661));
U_F10662: entity F port map(lamdaA => P(10)(662),lamdaB => P(10)(663),lamdaOut => P(9)(662));
U_G10663: entity G port map(lamdaA => P(10)(662),lamdaB => P(10)(663),s => s(10)(331),lamdaOut => P(9)(663));
U_F10664: entity F port map(lamdaA => P(10)(664),lamdaB => P(10)(665),lamdaOut => P(9)(664));
U_G10665: entity G port map(lamdaA => P(10)(664),lamdaB => P(10)(665),s => s(10)(332),lamdaOut => P(9)(665));
U_F10666: entity F port map(lamdaA => P(10)(666),lamdaB => P(10)(667),lamdaOut => P(9)(666));
U_G10667: entity G port map(lamdaA => P(10)(666),lamdaB => P(10)(667),s => s(10)(333),lamdaOut => P(9)(667));
U_F10668: entity F port map(lamdaA => P(10)(668),lamdaB => P(10)(669),lamdaOut => P(9)(668));
U_G10669: entity G port map(lamdaA => P(10)(668),lamdaB => P(10)(669),s => s(10)(334),lamdaOut => P(9)(669));
U_F10670: entity F port map(lamdaA => P(10)(670),lamdaB => P(10)(671),lamdaOut => P(9)(670));
U_G10671: entity G port map(lamdaA => P(10)(670),lamdaB => P(10)(671),s => s(10)(335),lamdaOut => P(9)(671));
U_F10672: entity F port map(lamdaA => P(10)(672),lamdaB => P(10)(673),lamdaOut => P(9)(672));
U_G10673: entity G port map(lamdaA => P(10)(672),lamdaB => P(10)(673),s => s(10)(336),lamdaOut => P(9)(673));
U_F10674: entity F port map(lamdaA => P(10)(674),lamdaB => P(10)(675),lamdaOut => P(9)(674));
U_G10675: entity G port map(lamdaA => P(10)(674),lamdaB => P(10)(675),s => s(10)(337),lamdaOut => P(9)(675));
U_F10676: entity F port map(lamdaA => P(10)(676),lamdaB => P(10)(677),lamdaOut => P(9)(676));
U_G10677: entity G port map(lamdaA => P(10)(676),lamdaB => P(10)(677),s => s(10)(338),lamdaOut => P(9)(677));
U_F10678: entity F port map(lamdaA => P(10)(678),lamdaB => P(10)(679),lamdaOut => P(9)(678));
U_G10679: entity G port map(lamdaA => P(10)(678),lamdaB => P(10)(679),s => s(10)(339),lamdaOut => P(9)(679));
U_F10680: entity F port map(lamdaA => P(10)(680),lamdaB => P(10)(681),lamdaOut => P(9)(680));
U_G10681: entity G port map(lamdaA => P(10)(680),lamdaB => P(10)(681),s => s(10)(340),lamdaOut => P(9)(681));
U_F10682: entity F port map(lamdaA => P(10)(682),lamdaB => P(10)(683),lamdaOut => P(9)(682));
U_G10683: entity G port map(lamdaA => P(10)(682),lamdaB => P(10)(683),s => s(10)(341),lamdaOut => P(9)(683));
U_F10684: entity F port map(lamdaA => P(10)(684),lamdaB => P(10)(685),lamdaOut => P(9)(684));
U_G10685: entity G port map(lamdaA => P(10)(684),lamdaB => P(10)(685),s => s(10)(342),lamdaOut => P(9)(685));
U_F10686: entity F port map(lamdaA => P(10)(686),lamdaB => P(10)(687),lamdaOut => P(9)(686));
U_G10687: entity G port map(lamdaA => P(10)(686),lamdaB => P(10)(687),s => s(10)(343),lamdaOut => P(9)(687));
U_F10688: entity F port map(lamdaA => P(10)(688),lamdaB => P(10)(689),lamdaOut => P(9)(688));
U_G10689: entity G port map(lamdaA => P(10)(688),lamdaB => P(10)(689),s => s(10)(344),lamdaOut => P(9)(689));
U_F10690: entity F port map(lamdaA => P(10)(690),lamdaB => P(10)(691),lamdaOut => P(9)(690));
U_G10691: entity G port map(lamdaA => P(10)(690),lamdaB => P(10)(691),s => s(10)(345),lamdaOut => P(9)(691));
U_F10692: entity F port map(lamdaA => P(10)(692),lamdaB => P(10)(693),lamdaOut => P(9)(692));
U_G10693: entity G port map(lamdaA => P(10)(692),lamdaB => P(10)(693),s => s(10)(346),lamdaOut => P(9)(693));
U_F10694: entity F port map(lamdaA => P(10)(694),lamdaB => P(10)(695),lamdaOut => P(9)(694));
U_G10695: entity G port map(lamdaA => P(10)(694),lamdaB => P(10)(695),s => s(10)(347),lamdaOut => P(9)(695));
U_F10696: entity F port map(lamdaA => P(10)(696),lamdaB => P(10)(697),lamdaOut => P(9)(696));
U_G10697: entity G port map(lamdaA => P(10)(696),lamdaB => P(10)(697),s => s(10)(348),lamdaOut => P(9)(697));
U_F10698: entity F port map(lamdaA => P(10)(698),lamdaB => P(10)(699),lamdaOut => P(9)(698));
U_G10699: entity G port map(lamdaA => P(10)(698),lamdaB => P(10)(699),s => s(10)(349),lamdaOut => P(9)(699));
U_F10700: entity F port map(lamdaA => P(10)(700),lamdaB => P(10)(701),lamdaOut => P(9)(700));
U_G10701: entity G port map(lamdaA => P(10)(700),lamdaB => P(10)(701),s => s(10)(350),lamdaOut => P(9)(701));
U_F10702: entity F port map(lamdaA => P(10)(702),lamdaB => P(10)(703),lamdaOut => P(9)(702));
U_G10703: entity G port map(lamdaA => P(10)(702),lamdaB => P(10)(703),s => s(10)(351),lamdaOut => P(9)(703));
U_F10704: entity F port map(lamdaA => P(10)(704),lamdaB => P(10)(705),lamdaOut => P(9)(704));
U_G10705: entity G port map(lamdaA => P(10)(704),lamdaB => P(10)(705),s => s(10)(352),lamdaOut => P(9)(705));
U_F10706: entity F port map(lamdaA => P(10)(706),lamdaB => P(10)(707),lamdaOut => P(9)(706));
U_G10707: entity G port map(lamdaA => P(10)(706),lamdaB => P(10)(707),s => s(10)(353),lamdaOut => P(9)(707));
U_F10708: entity F port map(lamdaA => P(10)(708),lamdaB => P(10)(709),lamdaOut => P(9)(708));
U_G10709: entity G port map(lamdaA => P(10)(708),lamdaB => P(10)(709),s => s(10)(354),lamdaOut => P(9)(709));
U_F10710: entity F port map(lamdaA => P(10)(710),lamdaB => P(10)(711),lamdaOut => P(9)(710));
U_G10711: entity G port map(lamdaA => P(10)(710),lamdaB => P(10)(711),s => s(10)(355),lamdaOut => P(9)(711));
U_F10712: entity F port map(lamdaA => P(10)(712),lamdaB => P(10)(713),lamdaOut => P(9)(712));
U_G10713: entity G port map(lamdaA => P(10)(712),lamdaB => P(10)(713),s => s(10)(356),lamdaOut => P(9)(713));
U_F10714: entity F port map(lamdaA => P(10)(714),lamdaB => P(10)(715),lamdaOut => P(9)(714));
U_G10715: entity G port map(lamdaA => P(10)(714),lamdaB => P(10)(715),s => s(10)(357),lamdaOut => P(9)(715));
U_F10716: entity F port map(lamdaA => P(10)(716),lamdaB => P(10)(717),lamdaOut => P(9)(716));
U_G10717: entity G port map(lamdaA => P(10)(716),lamdaB => P(10)(717),s => s(10)(358),lamdaOut => P(9)(717));
U_F10718: entity F port map(lamdaA => P(10)(718),lamdaB => P(10)(719),lamdaOut => P(9)(718));
U_G10719: entity G port map(lamdaA => P(10)(718),lamdaB => P(10)(719),s => s(10)(359),lamdaOut => P(9)(719));
U_F10720: entity F port map(lamdaA => P(10)(720),lamdaB => P(10)(721),lamdaOut => P(9)(720));
U_G10721: entity G port map(lamdaA => P(10)(720),lamdaB => P(10)(721),s => s(10)(360),lamdaOut => P(9)(721));
U_F10722: entity F port map(lamdaA => P(10)(722),lamdaB => P(10)(723),lamdaOut => P(9)(722));
U_G10723: entity G port map(lamdaA => P(10)(722),lamdaB => P(10)(723),s => s(10)(361),lamdaOut => P(9)(723));
U_F10724: entity F port map(lamdaA => P(10)(724),lamdaB => P(10)(725),lamdaOut => P(9)(724));
U_G10725: entity G port map(lamdaA => P(10)(724),lamdaB => P(10)(725),s => s(10)(362),lamdaOut => P(9)(725));
U_F10726: entity F port map(lamdaA => P(10)(726),lamdaB => P(10)(727),lamdaOut => P(9)(726));
U_G10727: entity G port map(lamdaA => P(10)(726),lamdaB => P(10)(727),s => s(10)(363),lamdaOut => P(9)(727));
U_F10728: entity F port map(lamdaA => P(10)(728),lamdaB => P(10)(729),lamdaOut => P(9)(728));
U_G10729: entity G port map(lamdaA => P(10)(728),lamdaB => P(10)(729),s => s(10)(364),lamdaOut => P(9)(729));
U_F10730: entity F port map(lamdaA => P(10)(730),lamdaB => P(10)(731),lamdaOut => P(9)(730));
U_G10731: entity G port map(lamdaA => P(10)(730),lamdaB => P(10)(731),s => s(10)(365),lamdaOut => P(9)(731));
U_F10732: entity F port map(lamdaA => P(10)(732),lamdaB => P(10)(733),lamdaOut => P(9)(732));
U_G10733: entity G port map(lamdaA => P(10)(732),lamdaB => P(10)(733),s => s(10)(366),lamdaOut => P(9)(733));
U_F10734: entity F port map(lamdaA => P(10)(734),lamdaB => P(10)(735),lamdaOut => P(9)(734));
U_G10735: entity G port map(lamdaA => P(10)(734),lamdaB => P(10)(735),s => s(10)(367),lamdaOut => P(9)(735));
U_F10736: entity F port map(lamdaA => P(10)(736),lamdaB => P(10)(737),lamdaOut => P(9)(736));
U_G10737: entity G port map(lamdaA => P(10)(736),lamdaB => P(10)(737),s => s(10)(368),lamdaOut => P(9)(737));
U_F10738: entity F port map(lamdaA => P(10)(738),lamdaB => P(10)(739),lamdaOut => P(9)(738));
U_G10739: entity G port map(lamdaA => P(10)(738),lamdaB => P(10)(739),s => s(10)(369),lamdaOut => P(9)(739));
U_F10740: entity F port map(lamdaA => P(10)(740),lamdaB => P(10)(741),lamdaOut => P(9)(740));
U_G10741: entity G port map(lamdaA => P(10)(740),lamdaB => P(10)(741),s => s(10)(370),lamdaOut => P(9)(741));
U_F10742: entity F port map(lamdaA => P(10)(742),lamdaB => P(10)(743),lamdaOut => P(9)(742));
U_G10743: entity G port map(lamdaA => P(10)(742),lamdaB => P(10)(743),s => s(10)(371),lamdaOut => P(9)(743));
U_F10744: entity F port map(lamdaA => P(10)(744),lamdaB => P(10)(745),lamdaOut => P(9)(744));
U_G10745: entity G port map(lamdaA => P(10)(744),lamdaB => P(10)(745),s => s(10)(372),lamdaOut => P(9)(745));
U_F10746: entity F port map(lamdaA => P(10)(746),lamdaB => P(10)(747),lamdaOut => P(9)(746));
U_G10747: entity G port map(lamdaA => P(10)(746),lamdaB => P(10)(747),s => s(10)(373),lamdaOut => P(9)(747));
U_F10748: entity F port map(lamdaA => P(10)(748),lamdaB => P(10)(749),lamdaOut => P(9)(748));
U_G10749: entity G port map(lamdaA => P(10)(748),lamdaB => P(10)(749),s => s(10)(374),lamdaOut => P(9)(749));
U_F10750: entity F port map(lamdaA => P(10)(750),lamdaB => P(10)(751),lamdaOut => P(9)(750));
U_G10751: entity G port map(lamdaA => P(10)(750),lamdaB => P(10)(751),s => s(10)(375),lamdaOut => P(9)(751));
U_F10752: entity F port map(lamdaA => P(10)(752),lamdaB => P(10)(753),lamdaOut => P(9)(752));
U_G10753: entity G port map(lamdaA => P(10)(752),lamdaB => P(10)(753),s => s(10)(376),lamdaOut => P(9)(753));
U_F10754: entity F port map(lamdaA => P(10)(754),lamdaB => P(10)(755),lamdaOut => P(9)(754));
U_G10755: entity G port map(lamdaA => P(10)(754),lamdaB => P(10)(755),s => s(10)(377),lamdaOut => P(9)(755));
U_F10756: entity F port map(lamdaA => P(10)(756),lamdaB => P(10)(757),lamdaOut => P(9)(756));
U_G10757: entity G port map(lamdaA => P(10)(756),lamdaB => P(10)(757),s => s(10)(378),lamdaOut => P(9)(757));
U_F10758: entity F port map(lamdaA => P(10)(758),lamdaB => P(10)(759),lamdaOut => P(9)(758));
U_G10759: entity G port map(lamdaA => P(10)(758),lamdaB => P(10)(759),s => s(10)(379),lamdaOut => P(9)(759));
U_F10760: entity F port map(lamdaA => P(10)(760),lamdaB => P(10)(761),lamdaOut => P(9)(760));
U_G10761: entity G port map(lamdaA => P(10)(760),lamdaB => P(10)(761),s => s(10)(380),lamdaOut => P(9)(761));
U_F10762: entity F port map(lamdaA => P(10)(762),lamdaB => P(10)(763),lamdaOut => P(9)(762));
U_G10763: entity G port map(lamdaA => P(10)(762),lamdaB => P(10)(763),s => s(10)(381),lamdaOut => P(9)(763));
U_F10764: entity F port map(lamdaA => P(10)(764),lamdaB => P(10)(765),lamdaOut => P(9)(764));
U_G10765: entity G port map(lamdaA => P(10)(764),lamdaB => P(10)(765),s => s(10)(382),lamdaOut => P(9)(765));
U_F10766: entity F port map(lamdaA => P(10)(766),lamdaB => P(10)(767),lamdaOut => P(9)(766));
U_G10767: entity G port map(lamdaA => P(10)(766),lamdaB => P(10)(767),s => s(10)(383),lamdaOut => P(9)(767));
U_F10768: entity F port map(lamdaA => P(10)(768),lamdaB => P(10)(769),lamdaOut => P(9)(768));
U_G10769: entity G port map(lamdaA => P(10)(768),lamdaB => P(10)(769),s => s(10)(384),lamdaOut => P(9)(769));
U_F10770: entity F port map(lamdaA => P(10)(770),lamdaB => P(10)(771),lamdaOut => P(9)(770));
U_G10771: entity G port map(lamdaA => P(10)(770),lamdaB => P(10)(771),s => s(10)(385),lamdaOut => P(9)(771));
U_F10772: entity F port map(lamdaA => P(10)(772),lamdaB => P(10)(773),lamdaOut => P(9)(772));
U_G10773: entity G port map(lamdaA => P(10)(772),lamdaB => P(10)(773),s => s(10)(386),lamdaOut => P(9)(773));
U_F10774: entity F port map(lamdaA => P(10)(774),lamdaB => P(10)(775),lamdaOut => P(9)(774));
U_G10775: entity G port map(lamdaA => P(10)(774),lamdaB => P(10)(775),s => s(10)(387),lamdaOut => P(9)(775));
U_F10776: entity F port map(lamdaA => P(10)(776),lamdaB => P(10)(777),lamdaOut => P(9)(776));
U_G10777: entity G port map(lamdaA => P(10)(776),lamdaB => P(10)(777),s => s(10)(388),lamdaOut => P(9)(777));
U_F10778: entity F port map(lamdaA => P(10)(778),lamdaB => P(10)(779),lamdaOut => P(9)(778));
U_G10779: entity G port map(lamdaA => P(10)(778),lamdaB => P(10)(779),s => s(10)(389),lamdaOut => P(9)(779));
U_F10780: entity F port map(lamdaA => P(10)(780),lamdaB => P(10)(781),lamdaOut => P(9)(780));
U_G10781: entity G port map(lamdaA => P(10)(780),lamdaB => P(10)(781),s => s(10)(390),lamdaOut => P(9)(781));
U_F10782: entity F port map(lamdaA => P(10)(782),lamdaB => P(10)(783),lamdaOut => P(9)(782));
U_G10783: entity G port map(lamdaA => P(10)(782),lamdaB => P(10)(783),s => s(10)(391),lamdaOut => P(9)(783));
U_F10784: entity F port map(lamdaA => P(10)(784),lamdaB => P(10)(785),lamdaOut => P(9)(784));
U_G10785: entity G port map(lamdaA => P(10)(784),lamdaB => P(10)(785),s => s(10)(392),lamdaOut => P(9)(785));
U_F10786: entity F port map(lamdaA => P(10)(786),lamdaB => P(10)(787),lamdaOut => P(9)(786));
U_G10787: entity G port map(lamdaA => P(10)(786),lamdaB => P(10)(787),s => s(10)(393),lamdaOut => P(9)(787));
U_F10788: entity F port map(lamdaA => P(10)(788),lamdaB => P(10)(789),lamdaOut => P(9)(788));
U_G10789: entity G port map(lamdaA => P(10)(788),lamdaB => P(10)(789),s => s(10)(394),lamdaOut => P(9)(789));
U_F10790: entity F port map(lamdaA => P(10)(790),lamdaB => P(10)(791),lamdaOut => P(9)(790));
U_G10791: entity G port map(lamdaA => P(10)(790),lamdaB => P(10)(791),s => s(10)(395),lamdaOut => P(9)(791));
U_F10792: entity F port map(lamdaA => P(10)(792),lamdaB => P(10)(793),lamdaOut => P(9)(792));
U_G10793: entity G port map(lamdaA => P(10)(792),lamdaB => P(10)(793),s => s(10)(396),lamdaOut => P(9)(793));
U_F10794: entity F port map(lamdaA => P(10)(794),lamdaB => P(10)(795),lamdaOut => P(9)(794));
U_G10795: entity G port map(lamdaA => P(10)(794),lamdaB => P(10)(795),s => s(10)(397),lamdaOut => P(9)(795));
U_F10796: entity F port map(lamdaA => P(10)(796),lamdaB => P(10)(797),lamdaOut => P(9)(796));
U_G10797: entity G port map(lamdaA => P(10)(796),lamdaB => P(10)(797),s => s(10)(398),lamdaOut => P(9)(797));
U_F10798: entity F port map(lamdaA => P(10)(798),lamdaB => P(10)(799),lamdaOut => P(9)(798));
U_G10799: entity G port map(lamdaA => P(10)(798),lamdaB => P(10)(799),s => s(10)(399),lamdaOut => P(9)(799));
U_F10800: entity F port map(lamdaA => P(10)(800),lamdaB => P(10)(801),lamdaOut => P(9)(800));
U_G10801: entity G port map(lamdaA => P(10)(800),lamdaB => P(10)(801),s => s(10)(400),lamdaOut => P(9)(801));
U_F10802: entity F port map(lamdaA => P(10)(802),lamdaB => P(10)(803),lamdaOut => P(9)(802));
U_G10803: entity G port map(lamdaA => P(10)(802),lamdaB => P(10)(803),s => s(10)(401),lamdaOut => P(9)(803));
U_F10804: entity F port map(lamdaA => P(10)(804),lamdaB => P(10)(805),lamdaOut => P(9)(804));
U_G10805: entity G port map(lamdaA => P(10)(804),lamdaB => P(10)(805),s => s(10)(402),lamdaOut => P(9)(805));
U_F10806: entity F port map(lamdaA => P(10)(806),lamdaB => P(10)(807),lamdaOut => P(9)(806));
U_G10807: entity G port map(lamdaA => P(10)(806),lamdaB => P(10)(807),s => s(10)(403),lamdaOut => P(9)(807));
U_F10808: entity F port map(lamdaA => P(10)(808),lamdaB => P(10)(809),lamdaOut => P(9)(808));
U_G10809: entity G port map(lamdaA => P(10)(808),lamdaB => P(10)(809),s => s(10)(404),lamdaOut => P(9)(809));
U_F10810: entity F port map(lamdaA => P(10)(810),lamdaB => P(10)(811),lamdaOut => P(9)(810));
U_G10811: entity G port map(lamdaA => P(10)(810),lamdaB => P(10)(811),s => s(10)(405),lamdaOut => P(9)(811));
U_F10812: entity F port map(lamdaA => P(10)(812),lamdaB => P(10)(813),lamdaOut => P(9)(812));
U_G10813: entity G port map(lamdaA => P(10)(812),lamdaB => P(10)(813),s => s(10)(406),lamdaOut => P(9)(813));
U_F10814: entity F port map(lamdaA => P(10)(814),lamdaB => P(10)(815),lamdaOut => P(9)(814));
U_G10815: entity G port map(lamdaA => P(10)(814),lamdaB => P(10)(815),s => s(10)(407),lamdaOut => P(9)(815));
U_F10816: entity F port map(lamdaA => P(10)(816),lamdaB => P(10)(817),lamdaOut => P(9)(816));
U_G10817: entity G port map(lamdaA => P(10)(816),lamdaB => P(10)(817),s => s(10)(408),lamdaOut => P(9)(817));
U_F10818: entity F port map(lamdaA => P(10)(818),lamdaB => P(10)(819),lamdaOut => P(9)(818));
U_G10819: entity G port map(lamdaA => P(10)(818),lamdaB => P(10)(819),s => s(10)(409),lamdaOut => P(9)(819));
U_F10820: entity F port map(lamdaA => P(10)(820),lamdaB => P(10)(821),lamdaOut => P(9)(820));
U_G10821: entity G port map(lamdaA => P(10)(820),lamdaB => P(10)(821),s => s(10)(410),lamdaOut => P(9)(821));
U_F10822: entity F port map(lamdaA => P(10)(822),lamdaB => P(10)(823),lamdaOut => P(9)(822));
U_G10823: entity G port map(lamdaA => P(10)(822),lamdaB => P(10)(823),s => s(10)(411),lamdaOut => P(9)(823));
U_F10824: entity F port map(lamdaA => P(10)(824),lamdaB => P(10)(825),lamdaOut => P(9)(824));
U_G10825: entity G port map(lamdaA => P(10)(824),lamdaB => P(10)(825),s => s(10)(412),lamdaOut => P(9)(825));
U_F10826: entity F port map(lamdaA => P(10)(826),lamdaB => P(10)(827),lamdaOut => P(9)(826));
U_G10827: entity G port map(lamdaA => P(10)(826),lamdaB => P(10)(827),s => s(10)(413),lamdaOut => P(9)(827));
U_F10828: entity F port map(lamdaA => P(10)(828),lamdaB => P(10)(829),lamdaOut => P(9)(828));
U_G10829: entity G port map(lamdaA => P(10)(828),lamdaB => P(10)(829),s => s(10)(414),lamdaOut => P(9)(829));
U_F10830: entity F port map(lamdaA => P(10)(830),lamdaB => P(10)(831),lamdaOut => P(9)(830));
U_G10831: entity G port map(lamdaA => P(10)(830),lamdaB => P(10)(831),s => s(10)(415),lamdaOut => P(9)(831));
U_F10832: entity F port map(lamdaA => P(10)(832),lamdaB => P(10)(833),lamdaOut => P(9)(832));
U_G10833: entity G port map(lamdaA => P(10)(832),lamdaB => P(10)(833),s => s(10)(416),lamdaOut => P(9)(833));
U_F10834: entity F port map(lamdaA => P(10)(834),lamdaB => P(10)(835),lamdaOut => P(9)(834));
U_G10835: entity G port map(lamdaA => P(10)(834),lamdaB => P(10)(835),s => s(10)(417),lamdaOut => P(9)(835));
U_F10836: entity F port map(lamdaA => P(10)(836),lamdaB => P(10)(837),lamdaOut => P(9)(836));
U_G10837: entity G port map(lamdaA => P(10)(836),lamdaB => P(10)(837),s => s(10)(418),lamdaOut => P(9)(837));
U_F10838: entity F port map(lamdaA => P(10)(838),lamdaB => P(10)(839),lamdaOut => P(9)(838));
U_G10839: entity G port map(lamdaA => P(10)(838),lamdaB => P(10)(839),s => s(10)(419),lamdaOut => P(9)(839));
U_F10840: entity F port map(lamdaA => P(10)(840),lamdaB => P(10)(841),lamdaOut => P(9)(840));
U_G10841: entity G port map(lamdaA => P(10)(840),lamdaB => P(10)(841),s => s(10)(420),lamdaOut => P(9)(841));
U_F10842: entity F port map(lamdaA => P(10)(842),lamdaB => P(10)(843),lamdaOut => P(9)(842));
U_G10843: entity G port map(lamdaA => P(10)(842),lamdaB => P(10)(843),s => s(10)(421),lamdaOut => P(9)(843));
U_F10844: entity F port map(lamdaA => P(10)(844),lamdaB => P(10)(845),lamdaOut => P(9)(844));
U_G10845: entity G port map(lamdaA => P(10)(844),lamdaB => P(10)(845),s => s(10)(422),lamdaOut => P(9)(845));
U_F10846: entity F port map(lamdaA => P(10)(846),lamdaB => P(10)(847),lamdaOut => P(9)(846));
U_G10847: entity G port map(lamdaA => P(10)(846),lamdaB => P(10)(847),s => s(10)(423),lamdaOut => P(9)(847));
U_F10848: entity F port map(lamdaA => P(10)(848),lamdaB => P(10)(849),lamdaOut => P(9)(848));
U_G10849: entity G port map(lamdaA => P(10)(848),lamdaB => P(10)(849),s => s(10)(424),lamdaOut => P(9)(849));
U_F10850: entity F port map(lamdaA => P(10)(850),lamdaB => P(10)(851),lamdaOut => P(9)(850));
U_G10851: entity G port map(lamdaA => P(10)(850),lamdaB => P(10)(851),s => s(10)(425),lamdaOut => P(9)(851));
U_F10852: entity F port map(lamdaA => P(10)(852),lamdaB => P(10)(853),lamdaOut => P(9)(852));
U_G10853: entity G port map(lamdaA => P(10)(852),lamdaB => P(10)(853),s => s(10)(426),lamdaOut => P(9)(853));
U_F10854: entity F port map(lamdaA => P(10)(854),lamdaB => P(10)(855),lamdaOut => P(9)(854));
U_G10855: entity G port map(lamdaA => P(10)(854),lamdaB => P(10)(855),s => s(10)(427),lamdaOut => P(9)(855));
U_F10856: entity F port map(lamdaA => P(10)(856),lamdaB => P(10)(857),lamdaOut => P(9)(856));
U_G10857: entity G port map(lamdaA => P(10)(856),lamdaB => P(10)(857),s => s(10)(428),lamdaOut => P(9)(857));
U_F10858: entity F port map(lamdaA => P(10)(858),lamdaB => P(10)(859),lamdaOut => P(9)(858));
U_G10859: entity G port map(lamdaA => P(10)(858),lamdaB => P(10)(859),s => s(10)(429),lamdaOut => P(9)(859));
U_F10860: entity F port map(lamdaA => P(10)(860),lamdaB => P(10)(861),lamdaOut => P(9)(860));
U_G10861: entity G port map(lamdaA => P(10)(860),lamdaB => P(10)(861),s => s(10)(430),lamdaOut => P(9)(861));
U_F10862: entity F port map(lamdaA => P(10)(862),lamdaB => P(10)(863),lamdaOut => P(9)(862));
U_G10863: entity G port map(lamdaA => P(10)(862),lamdaB => P(10)(863),s => s(10)(431),lamdaOut => P(9)(863));
U_F10864: entity F port map(lamdaA => P(10)(864),lamdaB => P(10)(865),lamdaOut => P(9)(864));
U_G10865: entity G port map(lamdaA => P(10)(864),lamdaB => P(10)(865),s => s(10)(432),lamdaOut => P(9)(865));
U_F10866: entity F port map(lamdaA => P(10)(866),lamdaB => P(10)(867),lamdaOut => P(9)(866));
U_G10867: entity G port map(lamdaA => P(10)(866),lamdaB => P(10)(867),s => s(10)(433),lamdaOut => P(9)(867));
U_F10868: entity F port map(lamdaA => P(10)(868),lamdaB => P(10)(869),lamdaOut => P(9)(868));
U_G10869: entity G port map(lamdaA => P(10)(868),lamdaB => P(10)(869),s => s(10)(434),lamdaOut => P(9)(869));
U_F10870: entity F port map(lamdaA => P(10)(870),lamdaB => P(10)(871),lamdaOut => P(9)(870));
U_G10871: entity G port map(lamdaA => P(10)(870),lamdaB => P(10)(871),s => s(10)(435),lamdaOut => P(9)(871));
U_F10872: entity F port map(lamdaA => P(10)(872),lamdaB => P(10)(873),lamdaOut => P(9)(872));
U_G10873: entity G port map(lamdaA => P(10)(872),lamdaB => P(10)(873),s => s(10)(436),lamdaOut => P(9)(873));
U_F10874: entity F port map(lamdaA => P(10)(874),lamdaB => P(10)(875),lamdaOut => P(9)(874));
U_G10875: entity G port map(lamdaA => P(10)(874),lamdaB => P(10)(875),s => s(10)(437),lamdaOut => P(9)(875));
U_F10876: entity F port map(lamdaA => P(10)(876),lamdaB => P(10)(877),lamdaOut => P(9)(876));
U_G10877: entity G port map(lamdaA => P(10)(876),lamdaB => P(10)(877),s => s(10)(438),lamdaOut => P(9)(877));
U_F10878: entity F port map(lamdaA => P(10)(878),lamdaB => P(10)(879),lamdaOut => P(9)(878));
U_G10879: entity G port map(lamdaA => P(10)(878),lamdaB => P(10)(879),s => s(10)(439),lamdaOut => P(9)(879));
U_F10880: entity F port map(lamdaA => P(10)(880),lamdaB => P(10)(881),lamdaOut => P(9)(880));
U_G10881: entity G port map(lamdaA => P(10)(880),lamdaB => P(10)(881),s => s(10)(440),lamdaOut => P(9)(881));
U_F10882: entity F port map(lamdaA => P(10)(882),lamdaB => P(10)(883),lamdaOut => P(9)(882));
U_G10883: entity G port map(lamdaA => P(10)(882),lamdaB => P(10)(883),s => s(10)(441),lamdaOut => P(9)(883));
U_F10884: entity F port map(lamdaA => P(10)(884),lamdaB => P(10)(885),lamdaOut => P(9)(884));
U_G10885: entity G port map(lamdaA => P(10)(884),lamdaB => P(10)(885),s => s(10)(442),lamdaOut => P(9)(885));
U_F10886: entity F port map(lamdaA => P(10)(886),lamdaB => P(10)(887),lamdaOut => P(9)(886));
U_G10887: entity G port map(lamdaA => P(10)(886),lamdaB => P(10)(887),s => s(10)(443),lamdaOut => P(9)(887));
U_F10888: entity F port map(lamdaA => P(10)(888),lamdaB => P(10)(889),lamdaOut => P(9)(888));
U_G10889: entity G port map(lamdaA => P(10)(888),lamdaB => P(10)(889),s => s(10)(444),lamdaOut => P(9)(889));
U_F10890: entity F port map(lamdaA => P(10)(890),lamdaB => P(10)(891),lamdaOut => P(9)(890));
U_G10891: entity G port map(lamdaA => P(10)(890),lamdaB => P(10)(891),s => s(10)(445),lamdaOut => P(9)(891));
U_F10892: entity F port map(lamdaA => P(10)(892),lamdaB => P(10)(893),lamdaOut => P(9)(892));
U_G10893: entity G port map(lamdaA => P(10)(892),lamdaB => P(10)(893),s => s(10)(446),lamdaOut => P(9)(893));
U_F10894: entity F port map(lamdaA => P(10)(894),lamdaB => P(10)(895),lamdaOut => P(9)(894));
U_G10895: entity G port map(lamdaA => P(10)(894),lamdaB => P(10)(895),s => s(10)(447),lamdaOut => P(9)(895));
U_F10896: entity F port map(lamdaA => P(10)(896),lamdaB => P(10)(897),lamdaOut => P(9)(896));
U_G10897: entity G port map(lamdaA => P(10)(896),lamdaB => P(10)(897),s => s(10)(448),lamdaOut => P(9)(897));
U_F10898: entity F port map(lamdaA => P(10)(898),lamdaB => P(10)(899),lamdaOut => P(9)(898));
U_G10899: entity G port map(lamdaA => P(10)(898),lamdaB => P(10)(899),s => s(10)(449),lamdaOut => P(9)(899));
U_F10900: entity F port map(lamdaA => P(10)(900),lamdaB => P(10)(901),lamdaOut => P(9)(900));
U_G10901: entity G port map(lamdaA => P(10)(900),lamdaB => P(10)(901),s => s(10)(450),lamdaOut => P(9)(901));
U_F10902: entity F port map(lamdaA => P(10)(902),lamdaB => P(10)(903),lamdaOut => P(9)(902));
U_G10903: entity G port map(lamdaA => P(10)(902),lamdaB => P(10)(903),s => s(10)(451),lamdaOut => P(9)(903));
U_F10904: entity F port map(lamdaA => P(10)(904),lamdaB => P(10)(905),lamdaOut => P(9)(904));
U_G10905: entity G port map(lamdaA => P(10)(904),lamdaB => P(10)(905),s => s(10)(452),lamdaOut => P(9)(905));
U_F10906: entity F port map(lamdaA => P(10)(906),lamdaB => P(10)(907),lamdaOut => P(9)(906));
U_G10907: entity G port map(lamdaA => P(10)(906),lamdaB => P(10)(907),s => s(10)(453),lamdaOut => P(9)(907));
U_F10908: entity F port map(lamdaA => P(10)(908),lamdaB => P(10)(909),lamdaOut => P(9)(908));
U_G10909: entity G port map(lamdaA => P(10)(908),lamdaB => P(10)(909),s => s(10)(454),lamdaOut => P(9)(909));
U_F10910: entity F port map(lamdaA => P(10)(910),lamdaB => P(10)(911),lamdaOut => P(9)(910));
U_G10911: entity G port map(lamdaA => P(10)(910),lamdaB => P(10)(911),s => s(10)(455),lamdaOut => P(9)(911));
U_F10912: entity F port map(lamdaA => P(10)(912),lamdaB => P(10)(913),lamdaOut => P(9)(912));
U_G10913: entity G port map(lamdaA => P(10)(912),lamdaB => P(10)(913),s => s(10)(456),lamdaOut => P(9)(913));
U_F10914: entity F port map(lamdaA => P(10)(914),lamdaB => P(10)(915),lamdaOut => P(9)(914));
U_G10915: entity G port map(lamdaA => P(10)(914),lamdaB => P(10)(915),s => s(10)(457),lamdaOut => P(9)(915));
U_F10916: entity F port map(lamdaA => P(10)(916),lamdaB => P(10)(917),lamdaOut => P(9)(916));
U_G10917: entity G port map(lamdaA => P(10)(916),lamdaB => P(10)(917),s => s(10)(458),lamdaOut => P(9)(917));
U_F10918: entity F port map(lamdaA => P(10)(918),lamdaB => P(10)(919),lamdaOut => P(9)(918));
U_G10919: entity G port map(lamdaA => P(10)(918),lamdaB => P(10)(919),s => s(10)(459),lamdaOut => P(9)(919));
U_F10920: entity F port map(lamdaA => P(10)(920),lamdaB => P(10)(921),lamdaOut => P(9)(920));
U_G10921: entity G port map(lamdaA => P(10)(920),lamdaB => P(10)(921),s => s(10)(460),lamdaOut => P(9)(921));
U_F10922: entity F port map(lamdaA => P(10)(922),lamdaB => P(10)(923),lamdaOut => P(9)(922));
U_G10923: entity G port map(lamdaA => P(10)(922),lamdaB => P(10)(923),s => s(10)(461),lamdaOut => P(9)(923));
U_F10924: entity F port map(lamdaA => P(10)(924),lamdaB => P(10)(925),lamdaOut => P(9)(924));
U_G10925: entity G port map(lamdaA => P(10)(924),lamdaB => P(10)(925),s => s(10)(462),lamdaOut => P(9)(925));
U_F10926: entity F port map(lamdaA => P(10)(926),lamdaB => P(10)(927),lamdaOut => P(9)(926));
U_G10927: entity G port map(lamdaA => P(10)(926),lamdaB => P(10)(927),s => s(10)(463),lamdaOut => P(9)(927));
U_F10928: entity F port map(lamdaA => P(10)(928),lamdaB => P(10)(929),lamdaOut => P(9)(928));
U_G10929: entity G port map(lamdaA => P(10)(928),lamdaB => P(10)(929),s => s(10)(464),lamdaOut => P(9)(929));
U_F10930: entity F port map(lamdaA => P(10)(930),lamdaB => P(10)(931),lamdaOut => P(9)(930));
U_G10931: entity G port map(lamdaA => P(10)(930),lamdaB => P(10)(931),s => s(10)(465),lamdaOut => P(9)(931));
U_F10932: entity F port map(lamdaA => P(10)(932),lamdaB => P(10)(933),lamdaOut => P(9)(932));
U_G10933: entity G port map(lamdaA => P(10)(932),lamdaB => P(10)(933),s => s(10)(466),lamdaOut => P(9)(933));
U_F10934: entity F port map(lamdaA => P(10)(934),lamdaB => P(10)(935),lamdaOut => P(9)(934));
U_G10935: entity G port map(lamdaA => P(10)(934),lamdaB => P(10)(935),s => s(10)(467),lamdaOut => P(9)(935));
U_F10936: entity F port map(lamdaA => P(10)(936),lamdaB => P(10)(937),lamdaOut => P(9)(936));
U_G10937: entity G port map(lamdaA => P(10)(936),lamdaB => P(10)(937),s => s(10)(468),lamdaOut => P(9)(937));
U_F10938: entity F port map(lamdaA => P(10)(938),lamdaB => P(10)(939),lamdaOut => P(9)(938));
U_G10939: entity G port map(lamdaA => P(10)(938),lamdaB => P(10)(939),s => s(10)(469),lamdaOut => P(9)(939));
U_F10940: entity F port map(lamdaA => P(10)(940),lamdaB => P(10)(941),lamdaOut => P(9)(940));
U_G10941: entity G port map(lamdaA => P(10)(940),lamdaB => P(10)(941),s => s(10)(470),lamdaOut => P(9)(941));
U_F10942: entity F port map(lamdaA => P(10)(942),lamdaB => P(10)(943),lamdaOut => P(9)(942));
U_G10943: entity G port map(lamdaA => P(10)(942),lamdaB => P(10)(943),s => s(10)(471),lamdaOut => P(9)(943));
U_F10944: entity F port map(lamdaA => P(10)(944),lamdaB => P(10)(945),lamdaOut => P(9)(944));
U_G10945: entity G port map(lamdaA => P(10)(944),lamdaB => P(10)(945),s => s(10)(472),lamdaOut => P(9)(945));
U_F10946: entity F port map(lamdaA => P(10)(946),lamdaB => P(10)(947),lamdaOut => P(9)(946));
U_G10947: entity G port map(lamdaA => P(10)(946),lamdaB => P(10)(947),s => s(10)(473),lamdaOut => P(9)(947));
U_F10948: entity F port map(lamdaA => P(10)(948),lamdaB => P(10)(949),lamdaOut => P(9)(948));
U_G10949: entity G port map(lamdaA => P(10)(948),lamdaB => P(10)(949),s => s(10)(474),lamdaOut => P(9)(949));
U_F10950: entity F port map(lamdaA => P(10)(950),lamdaB => P(10)(951),lamdaOut => P(9)(950));
U_G10951: entity G port map(lamdaA => P(10)(950),lamdaB => P(10)(951),s => s(10)(475),lamdaOut => P(9)(951));
U_F10952: entity F port map(lamdaA => P(10)(952),lamdaB => P(10)(953),lamdaOut => P(9)(952));
U_G10953: entity G port map(lamdaA => P(10)(952),lamdaB => P(10)(953),s => s(10)(476),lamdaOut => P(9)(953));
U_F10954: entity F port map(lamdaA => P(10)(954),lamdaB => P(10)(955),lamdaOut => P(9)(954));
U_G10955: entity G port map(lamdaA => P(10)(954),lamdaB => P(10)(955),s => s(10)(477),lamdaOut => P(9)(955));
U_F10956: entity F port map(lamdaA => P(10)(956),lamdaB => P(10)(957),lamdaOut => P(9)(956));
U_G10957: entity G port map(lamdaA => P(10)(956),lamdaB => P(10)(957),s => s(10)(478),lamdaOut => P(9)(957));
U_F10958: entity F port map(lamdaA => P(10)(958),lamdaB => P(10)(959),lamdaOut => P(9)(958));
U_G10959: entity G port map(lamdaA => P(10)(958),lamdaB => P(10)(959),s => s(10)(479),lamdaOut => P(9)(959));
U_F10960: entity F port map(lamdaA => P(10)(960),lamdaB => P(10)(961),lamdaOut => P(9)(960));
U_G10961: entity G port map(lamdaA => P(10)(960),lamdaB => P(10)(961),s => s(10)(480),lamdaOut => P(9)(961));
U_F10962: entity F port map(lamdaA => P(10)(962),lamdaB => P(10)(963),lamdaOut => P(9)(962));
U_G10963: entity G port map(lamdaA => P(10)(962),lamdaB => P(10)(963),s => s(10)(481),lamdaOut => P(9)(963));
U_F10964: entity F port map(lamdaA => P(10)(964),lamdaB => P(10)(965),lamdaOut => P(9)(964));
U_G10965: entity G port map(lamdaA => P(10)(964),lamdaB => P(10)(965),s => s(10)(482),lamdaOut => P(9)(965));
U_F10966: entity F port map(lamdaA => P(10)(966),lamdaB => P(10)(967),lamdaOut => P(9)(966));
U_G10967: entity G port map(lamdaA => P(10)(966),lamdaB => P(10)(967),s => s(10)(483),lamdaOut => P(9)(967));
U_F10968: entity F port map(lamdaA => P(10)(968),lamdaB => P(10)(969),lamdaOut => P(9)(968));
U_G10969: entity G port map(lamdaA => P(10)(968),lamdaB => P(10)(969),s => s(10)(484),lamdaOut => P(9)(969));
U_F10970: entity F port map(lamdaA => P(10)(970),lamdaB => P(10)(971),lamdaOut => P(9)(970));
U_G10971: entity G port map(lamdaA => P(10)(970),lamdaB => P(10)(971),s => s(10)(485),lamdaOut => P(9)(971));
U_F10972: entity F port map(lamdaA => P(10)(972),lamdaB => P(10)(973),lamdaOut => P(9)(972));
U_G10973: entity G port map(lamdaA => P(10)(972),lamdaB => P(10)(973),s => s(10)(486),lamdaOut => P(9)(973));
U_F10974: entity F port map(lamdaA => P(10)(974),lamdaB => P(10)(975),lamdaOut => P(9)(974));
U_G10975: entity G port map(lamdaA => P(10)(974),lamdaB => P(10)(975),s => s(10)(487),lamdaOut => P(9)(975));
U_F10976: entity F port map(lamdaA => P(10)(976),lamdaB => P(10)(977),lamdaOut => P(9)(976));
U_G10977: entity G port map(lamdaA => P(10)(976),lamdaB => P(10)(977),s => s(10)(488),lamdaOut => P(9)(977));
U_F10978: entity F port map(lamdaA => P(10)(978),lamdaB => P(10)(979),lamdaOut => P(9)(978));
U_G10979: entity G port map(lamdaA => P(10)(978),lamdaB => P(10)(979),s => s(10)(489),lamdaOut => P(9)(979));
U_F10980: entity F port map(lamdaA => P(10)(980),lamdaB => P(10)(981),lamdaOut => P(9)(980));
U_G10981: entity G port map(lamdaA => P(10)(980),lamdaB => P(10)(981),s => s(10)(490),lamdaOut => P(9)(981));
U_F10982: entity F port map(lamdaA => P(10)(982),lamdaB => P(10)(983),lamdaOut => P(9)(982));
U_G10983: entity G port map(lamdaA => P(10)(982),lamdaB => P(10)(983),s => s(10)(491),lamdaOut => P(9)(983));
U_F10984: entity F port map(lamdaA => P(10)(984),lamdaB => P(10)(985),lamdaOut => P(9)(984));
U_G10985: entity G port map(lamdaA => P(10)(984),lamdaB => P(10)(985),s => s(10)(492),lamdaOut => P(9)(985));
U_F10986: entity F port map(lamdaA => P(10)(986),lamdaB => P(10)(987),lamdaOut => P(9)(986));
U_G10987: entity G port map(lamdaA => P(10)(986),lamdaB => P(10)(987),s => s(10)(493),lamdaOut => P(9)(987));
U_F10988: entity F port map(lamdaA => P(10)(988),lamdaB => P(10)(989),lamdaOut => P(9)(988));
U_G10989: entity G port map(lamdaA => P(10)(988),lamdaB => P(10)(989),s => s(10)(494),lamdaOut => P(9)(989));
U_F10990: entity F port map(lamdaA => P(10)(990),lamdaB => P(10)(991),lamdaOut => P(9)(990));
U_G10991: entity G port map(lamdaA => P(10)(990),lamdaB => P(10)(991),s => s(10)(495),lamdaOut => P(9)(991));
U_F10992: entity F port map(lamdaA => P(10)(992),lamdaB => P(10)(993),lamdaOut => P(9)(992));
U_G10993: entity G port map(lamdaA => P(10)(992),lamdaB => P(10)(993),s => s(10)(496),lamdaOut => P(9)(993));
U_F10994: entity F port map(lamdaA => P(10)(994),lamdaB => P(10)(995),lamdaOut => P(9)(994));
U_G10995: entity G port map(lamdaA => P(10)(994),lamdaB => P(10)(995),s => s(10)(497),lamdaOut => P(9)(995));
U_F10996: entity F port map(lamdaA => P(10)(996),lamdaB => P(10)(997),lamdaOut => P(9)(996));
U_G10997: entity G port map(lamdaA => P(10)(996),lamdaB => P(10)(997),s => s(10)(498),lamdaOut => P(9)(997));
U_F10998: entity F port map(lamdaA => P(10)(998),lamdaB => P(10)(999),lamdaOut => P(9)(998));
U_G10999: entity G port map(lamdaA => P(10)(998),lamdaB => P(10)(999),s => s(10)(499),lamdaOut => P(9)(999));
U_F101000: entity F port map(lamdaA => P(10)(1000),lamdaB => P(10)(1001),lamdaOut => P(9)(1000));
U_G101001: entity G port map(lamdaA => P(10)(1000),lamdaB => P(10)(1001),s => s(10)(500),lamdaOut => P(9)(1001));
U_F101002: entity F port map(lamdaA => P(10)(1002),lamdaB => P(10)(1003),lamdaOut => P(9)(1002));
U_G101003: entity G port map(lamdaA => P(10)(1002),lamdaB => P(10)(1003),s => s(10)(501),lamdaOut => P(9)(1003));
U_F101004: entity F port map(lamdaA => P(10)(1004),lamdaB => P(10)(1005),lamdaOut => P(9)(1004));
U_G101005: entity G port map(lamdaA => P(10)(1004),lamdaB => P(10)(1005),s => s(10)(502),lamdaOut => P(9)(1005));
U_F101006: entity F port map(lamdaA => P(10)(1006),lamdaB => P(10)(1007),lamdaOut => P(9)(1006));
U_G101007: entity G port map(lamdaA => P(10)(1006),lamdaB => P(10)(1007),s => s(10)(503),lamdaOut => P(9)(1007));
U_F101008: entity F port map(lamdaA => P(10)(1008),lamdaB => P(10)(1009),lamdaOut => P(9)(1008));
U_G101009: entity G port map(lamdaA => P(10)(1008),lamdaB => P(10)(1009),s => s(10)(504),lamdaOut => P(9)(1009));
U_F101010: entity F port map(lamdaA => P(10)(1010),lamdaB => P(10)(1011),lamdaOut => P(9)(1010));
U_G101011: entity G port map(lamdaA => P(10)(1010),lamdaB => P(10)(1011),s => s(10)(505),lamdaOut => P(9)(1011));
U_F101012: entity F port map(lamdaA => P(10)(1012),lamdaB => P(10)(1013),lamdaOut => P(9)(1012));
U_G101013: entity G port map(lamdaA => P(10)(1012),lamdaB => P(10)(1013),s => s(10)(506),lamdaOut => P(9)(1013));
U_F101014: entity F port map(lamdaA => P(10)(1014),lamdaB => P(10)(1015),lamdaOut => P(9)(1014));
U_G101015: entity G port map(lamdaA => P(10)(1014),lamdaB => P(10)(1015),s => s(10)(507),lamdaOut => P(9)(1015));
U_F101016: entity F port map(lamdaA => P(10)(1016),lamdaB => P(10)(1017),lamdaOut => P(9)(1016));
U_G101017: entity G port map(lamdaA => P(10)(1016),lamdaB => P(10)(1017),s => s(10)(508),lamdaOut => P(9)(1017));
U_F101018: entity F port map(lamdaA => P(10)(1018),lamdaB => P(10)(1019),lamdaOut => P(9)(1018));
U_G101019: entity G port map(lamdaA => P(10)(1018),lamdaB => P(10)(1019),s => s(10)(509),lamdaOut => P(9)(1019));
U_F101020: entity F port map(lamdaA => P(10)(1020),lamdaB => P(10)(1021),lamdaOut => P(9)(1020));
U_G101021: entity G port map(lamdaA => P(10)(1020),lamdaB => P(10)(1021),s => s(10)(510),lamdaOut => P(9)(1021));
U_F101022: entity F port map(lamdaA => P(10)(1022),lamdaB => P(10)(1023),lamdaOut => P(9)(1022));
U_G101023: entity G port map(lamdaA => P(10)(1022),lamdaB => P(10)(1023),s => s(10)(511),lamdaOut => P(9)(1023));
-- STAGE 8
U_F90: entity F port map(lamdaA => P(9)(0),lamdaB => P(9)(2),lamdaOut => P(8)(0));
U_F91: entity F port map(lamdaA => P(9)(1),lamdaB => P(9)(3),lamdaOut => P(8)(1));
U_G92: entity G port map(lamdaA => P(9)(0),lamdaB => P(9)(2),s => s(9)(0),lamdaOut => P(8)(2));
U_G93: entity G port map(lamdaA => P(9)(1),lamdaB => P(9)(3),s => s(9)(1),lamdaOut => P(8)(3));
U_F94: entity F port map(lamdaA => P(9)(4),lamdaB => P(9)(6),lamdaOut => P(8)(4));
U_F95: entity F port map(lamdaA => P(9)(5),lamdaB => P(9)(7),lamdaOut => P(8)(5));
U_G96: entity G port map(lamdaA => P(9)(4),lamdaB => P(9)(6),s => s(9)(2),lamdaOut => P(8)(6));
U_G97: entity G port map(lamdaA => P(9)(5),lamdaB => P(9)(7),s => s(9)(3),lamdaOut => P(8)(7));
U_F98: entity F port map(lamdaA => P(9)(8),lamdaB => P(9)(10),lamdaOut => P(8)(8));
U_F99: entity F port map(lamdaA => P(9)(9),lamdaB => P(9)(11),lamdaOut => P(8)(9));
U_G910: entity G port map(lamdaA => P(9)(8),lamdaB => P(9)(10),s => s(9)(4),lamdaOut => P(8)(10));
U_G911: entity G port map(lamdaA => P(9)(9),lamdaB => P(9)(11),s => s(9)(5),lamdaOut => P(8)(11));
U_F912: entity F port map(lamdaA => P(9)(12),lamdaB => P(9)(14),lamdaOut => P(8)(12));
U_F913: entity F port map(lamdaA => P(9)(13),lamdaB => P(9)(15),lamdaOut => P(8)(13));
U_G914: entity G port map(lamdaA => P(9)(12),lamdaB => P(9)(14),s => s(9)(6),lamdaOut => P(8)(14));
U_G915: entity G port map(lamdaA => P(9)(13),lamdaB => P(9)(15),s => s(9)(7),lamdaOut => P(8)(15));
U_F916: entity F port map(lamdaA => P(9)(16),lamdaB => P(9)(18),lamdaOut => P(8)(16));
U_F917: entity F port map(lamdaA => P(9)(17),lamdaB => P(9)(19),lamdaOut => P(8)(17));
U_G918: entity G port map(lamdaA => P(9)(16),lamdaB => P(9)(18),s => s(9)(8),lamdaOut => P(8)(18));
U_G919: entity G port map(lamdaA => P(9)(17),lamdaB => P(9)(19),s => s(9)(9),lamdaOut => P(8)(19));
U_F920: entity F port map(lamdaA => P(9)(20),lamdaB => P(9)(22),lamdaOut => P(8)(20));
U_F921: entity F port map(lamdaA => P(9)(21),lamdaB => P(9)(23),lamdaOut => P(8)(21));
U_G922: entity G port map(lamdaA => P(9)(20),lamdaB => P(9)(22),s => s(9)(10),lamdaOut => P(8)(22));
U_G923: entity G port map(lamdaA => P(9)(21),lamdaB => P(9)(23),s => s(9)(11),lamdaOut => P(8)(23));
U_F924: entity F port map(lamdaA => P(9)(24),lamdaB => P(9)(26),lamdaOut => P(8)(24));
U_F925: entity F port map(lamdaA => P(9)(25),lamdaB => P(9)(27),lamdaOut => P(8)(25));
U_G926: entity G port map(lamdaA => P(9)(24),lamdaB => P(9)(26),s => s(9)(12),lamdaOut => P(8)(26));
U_G927: entity G port map(lamdaA => P(9)(25),lamdaB => P(9)(27),s => s(9)(13),lamdaOut => P(8)(27));
U_F928: entity F port map(lamdaA => P(9)(28),lamdaB => P(9)(30),lamdaOut => P(8)(28));
U_F929: entity F port map(lamdaA => P(9)(29),lamdaB => P(9)(31),lamdaOut => P(8)(29));
U_G930: entity G port map(lamdaA => P(9)(28),lamdaB => P(9)(30),s => s(9)(14),lamdaOut => P(8)(30));
U_G931: entity G port map(lamdaA => P(9)(29),lamdaB => P(9)(31),s => s(9)(15),lamdaOut => P(8)(31));
U_F932: entity F port map(lamdaA => P(9)(32),lamdaB => P(9)(34),lamdaOut => P(8)(32));
U_F933: entity F port map(lamdaA => P(9)(33),lamdaB => P(9)(35),lamdaOut => P(8)(33));
U_G934: entity G port map(lamdaA => P(9)(32),lamdaB => P(9)(34),s => s(9)(16),lamdaOut => P(8)(34));
U_G935: entity G port map(lamdaA => P(9)(33),lamdaB => P(9)(35),s => s(9)(17),lamdaOut => P(8)(35));
U_F936: entity F port map(lamdaA => P(9)(36),lamdaB => P(9)(38),lamdaOut => P(8)(36));
U_F937: entity F port map(lamdaA => P(9)(37),lamdaB => P(9)(39),lamdaOut => P(8)(37));
U_G938: entity G port map(lamdaA => P(9)(36),lamdaB => P(9)(38),s => s(9)(18),lamdaOut => P(8)(38));
U_G939: entity G port map(lamdaA => P(9)(37),lamdaB => P(9)(39),s => s(9)(19),lamdaOut => P(8)(39));
U_F940: entity F port map(lamdaA => P(9)(40),lamdaB => P(9)(42),lamdaOut => P(8)(40));
U_F941: entity F port map(lamdaA => P(9)(41),lamdaB => P(9)(43),lamdaOut => P(8)(41));
U_G942: entity G port map(lamdaA => P(9)(40),lamdaB => P(9)(42),s => s(9)(20),lamdaOut => P(8)(42));
U_G943: entity G port map(lamdaA => P(9)(41),lamdaB => P(9)(43),s => s(9)(21),lamdaOut => P(8)(43));
U_F944: entity F port map(lamdaA => P(9)(44),lamdaB => P(9)(46),lamdaOut => P(8)(44));
U_F945: entity F port map(lamdaA => P(9)(45),lamdaB => P(9)(47),lamdaOut => P(8)(45));
U_G946: entity G port map(lamdaA => P(9)(44),lamdaB => P(9)(46),s => s(9)(22),lamdaOut => P(8)(46));
U_G947: entity G port map(lamdaA => P(9)(45),lamdaB => P(9)(47),s => s(9)(23),lamdaOut => P(8)(47));
U_F948: entity F port map(lamdaA => P(9)(48),lamdaB => P(9)(50),lamdaOut => P(8)(48));
U_F949: entity F port map(lamdaA => P(9)(49),lamdaB => P(9)(51),lamdaOut => P(8)(49));
U_G950: entity G port map(lamdaA => P(9)(48),lamdaB => P(9)(50),s => s(9)(24),lamdaOut => P(8)(50));
U_G951: entity G port map(lamdaA => P(9)(49),lamdaB => P(9)(51),s => s(9)(25),lamdaOut => P(8)(51));
U_F952: entity F port map(lamdaA => P(9)(52),lamdaB => P(9)(54),lamdaOut => P(8)(52));
U_F953: entity F port map(lamdaA => P(9)(53),lamdaB => P(9)(55),lamdaOut => P(8)(53));
U_G954: entity G port map(lamdaA => P(9)(52),lamdaB => P(9)(54),s => s(9)(26),lamdaOut => P(8)(54));
U_G955: entity G port map(lamdaA => P(9)(53),lamdaB => P(9)(55),s => s(9)(27),lamdaOut => P(8)(55));
U_F956: entity F port map(lamdaA => P(9)(56),lamdaB => P(9)(58),lamdaOut => P(8)(56));
U_F957: entity F port map(lamdaA => P(9)(57),lamdaB => P(9)(59),lamdaOut => P(8)(57));
U_G958: entity G port map(lamdaA => P(9)(56),lamdaB => P(9)(58),s => s(9)(28),lamdaOut => P(8)(58));
U_G959: entity G port map(lamdaA => P(9)(57),lamdaB => P(9)(59),s => s(9)(29),lamdaOut => P(8)(59));
U_F960: entity F port map(lamdaA => P(9)(60),lamdaB => P(9)(62),lamdaOut => P(8)(60));
U_F961: entity F port map(lamdaA => P(9)(61),lamdaB => P(9)(63),lamdaOut => P(8)(61));
U_G962: entity G port map(lamdaA => P(9)(60),lamdaB => P(9)(62),s => s(9)(30),lamdaOut => P(8)(62));
U_G963: entity G port map(lamdaA => P(9)(61),lamdaB => P(9)(63),s => s(9)(31),lamdaOut => P(8)(63));
U_F964: entity F port map(lamdaA => P(9)(64),lamdaB => P(9)(66),lamdaOut => P(8)(64));
U_F965: entity F port map(lamdaA => P(9)(65),lamdaB => P(9)(67),lamdaOut => P(8)(65));
U_G966: entity G port map(lamdaA => P(9)(64),lamdaB => P(9)(66),s => s(9)(32),lamdaOut => P(8)(66));
U_G967: entity G port map(lamdaA => P(9)(65),lamdaB => P(9)(67),s => s(9)(33),lamdaOut => P(8)(67));
U_F968: entity F port map(lamdaA => P(9)(68),lamdaB => P(9)(70),lamdaOut => P(8)(68));
U_F969: entity F port map(lamdaA => P(9)(69),lamdaB => P(9)(71),lamdaOut => P(8)(69));
U_G970: entity G port map(lamdaA => P(9)(68),lamdaB => P(9)(70),s => s(9)(34),lamdaOut => P(8)(70));
U_G971: entity G port map(lamdaA => P(9)(69),lamdaB => P(9)(71),s => s(9)(35),lamdaOut => P(8)(71));
U_F972: entity F port map(lamdaA => P(9)(72),lamdaB => P(9)(74),lamdaOut => P(8)(72));
U_F973: entity F port map(lamdaA => P(9)(73),lamdaB => P(9)(75),lamdaOut => P(8)(73));
U_G974: entity G port map(lamdaA => P(9)(72),lamdaB => P(9)(74),s => s(9)(36),lamdaOut => P(8)(74));
U_G975: entity G port map(lamdaA => P(9)(73),lamdaB => P(9)(75),s => s(9)(37),lamdaOut => P(8)(75));
U_F976: entity F port map(lamdaA => P(9)(76),lamdaB => P(9)(78),lamdaOut => P(8)(76));
U_F977: entity F port map(lamdaA => P(9)(77),lamdaB => P(9)(79),lamdaOut => P(8)(77));
U_G978: entity G port map(lamdaA => P(9)(76),lamdaB => P(9)(78),s => s(9)(38),lamdaOut => P(8)(78));
U_G979: entity G port map(lamdaA => P(9)(77),lamdaB => P(9)(79),s => s(9)(39),lamdaOut => P(8)(79));
U_F980: entity F port map(lamdaA => P(9)(80),lamdaB => P(9)(82),lamdaOut => P(8)(80));
U_F981: entity F port map(lamdaA => P(9)(81),lamdaB => P(9)(83),lamdaOut => P(8)(81));
U_G982: entity G port map(lamdaA => P(9)(80),lamdaB => P(9)(82),s => s(9)(40),lamdaOut => P(8)(82));
U_G983: entity G port map(lamdaA => P(9)(81),lamdaB => P(9)(83),s => s(9)(41),lamdaOut => P(8)(83));
U_F984: entity F port map(lamdaA => P(9)(84),lamdaB => P(9)(86),lamdaOut => P(8)(84));
U_F985: entity F port map(lamdaA => P(9)(85),lamdaB => P(9)(87),lamdaOut => P(8)(85));
U_G986: entity G port map(lamdaA => P(9)(84),lamdaB => P(9)(86),s => s(9)(42),lamdaOut => P(8)(86));
U_G987: entity G port map(lamdaA => P(9)(85),lamdaB => P(9)(87),s => s(9)(43),lamdaOut => P(8)(87));
U_F988: entity F port map(lamdaA => P(9)(88),lamdaB => P(9)(90),lamdaOut => P(8)(88));
U_F989: entity F port map(lamdaA => P(9)(89),lamdaB => P(9)(91),lamdaOut => P(8)(89));
U_G990: entity G port map(lamdaA => P(9)(88),lamdaB => P(9)(90),s => s(9)(44),lamdaOut => P(8)(90));
U_G991: entity G port map(lamdaA => P(9)(89),lamdaB => P(9)(91),s => s(9)(45),lamdaOut => P(8)(91));
U_F992: entity F port map(lamdaA => P(9)(92),lamdaB => P(9)(94),lamdaOut => P(8)(92));
U_F993: entity F port map(lamdaA => P(9)(93),lamdaB => P(9)(95),lamdaOut => P(8)(93));
U_G994: entity G port map(lamdaA => P(9)(92),lamdaB => P(9)(94),s => s(9)(46),lamdaOut => P(8)(94));
U_G995: entity G port map(lamdaA => P(9)(93),lamdaB => P(9)(95),s => s(9)(47),lamdaOut => P(8)(95));
U_F996: entity F port map(lamdaA => P(9)(96),lamdaB => P(9)(98),lamdaOut => P(8)(96));
U_F997: entity F port map(lamdaA => P(9)(97),lamdaB => P(9)(99),lamdaOut => P(8)(97));
U_G998: entity G port map(lamdaA => P(9)(96),lamdaB => P(9)(98),s => s(9)(48),lamdaOut => P(8)(98));
U_G999: entity G port map(lamdaA => P(9)(97),lamdaB => P(9)(99),s => s(9)(49),lamdaOut => P(8)(99));
U_F9100: entity F port map(lamdaA => P(9)(100),lamdaB => P(9)(102),lamdaOut => P(8)(100));
U_F9101: entity F port map(lamdaA => P(9)(101),lamdaB => P(9)(103),lamdaOut => P(8)(101));
U_G9102: entity G port map(lamdaA => P(9)(100),lamdaB => P(9)(102),s => s(9)(50),lamdaOut => P(8)(102));
U_G9103: entity G port map(lamdaA => P(9)(101),lamdaB => P(9)(103),s => s(9)(51),lamdaOut => P(8)(103));
U_F9104: entity F port map(lamdaA => P(9)(104),lamdaB => P(9)(106),lamdaOut => P(8)(104));
U_F9105: entity F port map(lamdaA => P(9)(105),lamdaB => P(9)(107),lamdaOut => P(8)(105));
U_G9106: entity G port map(lamdaA => P(9)(104),lamdaB => P(9)(106),s => s(9)(52),lamdaOut => P(8)(106));
U_G9107: entity G port map(lamdaA => P(9)(105),lamdaB => P(9)(107),s => s(9)(53),lamdaOut => P(8)(107));
U_F9108: entity F port map(lamdaA => P(9)(108),lamdaB => P(9)(110),lamdaOut => P(8)(108));
U_F9109: entity F port map(lamdaA => P(9)(109),lamdaB => P(9)(111),lamdaOut => P(8)(109));
U_G9110: entity G port map(lamdaA => P(9)(108),lamdaB => P(9)(110),s => s(9)(54),lamdaOut => P(8)(110));
U_G9111: entity G port map(lamdaA => P(9)(109),lamdaB => P(9)(111),s => s(9)(55),lamdaOut => P(8)(111));
U_F9112: entity F port map(lamdaA => P(9)(112),lamdaB => P(9)(114),lamdaOut => P(8)(112));
U_F9113: entity F port map(lamdaA => P(9)(113),lamdaB => P(9)(115),lamdaOut => P(8)(113));
U_G9114: entity G port map(lamdaA => P(9)(112),lamdaB => P(9)(114),s => s(9)(56),lamdaOut => P(8)(114));
U_G9115: entity G port map(lamdaA => P(9)(113),lamdaB => P(9)(115),s => s(9)(57),lamdaOut => P(8)(115));
U_F9116: entity F port map(lamdaA => P(9)(116),lamdaB => P(9)(118),lamdaOut => P(8)(116));
U_F9117: entity F port map(lamdaA => P(9)(117),lamdaB => P(9)(119),lamdaOut => P(8)(117));
U_G9118: entity G port map(lamdaA => P(9)(116),lamdaB => P(9)(118),s => s(9)(58),lamdaOut => P(8)(118));
U_G9119: entity G port map(lamdaA => P(9)(117),lamdaB => P(9)(119),s => s(9)(59),lamdaOut => P(8)(119));
U_F9120: entity F port map(lamdaA => P(9)(120),lamdaB => P(9)(122),lamdaOut => P(8)(120));
U_F9121: entity F port map(lamdaA => P(9)(121),lamdaB => P(9)(123),lamdaOut => P(8)(121));
U_G9122: entity G port map(lamdaA => P(9)(120),lamdaB => P(9)(122),s => s(9)(60),lamdaOut => P(8)(122));
U_G9123: entity G port map(lamdaA => P(9)(121),lamdaB => P(9)(123),s => s(9)(61),lamdaOut => P(8)(123));
U_F9124: entity F port map(lamdaA => P(9)(124),lamdaB => P(9)(126),lamdaOut => P(8)(124));
U_F9125: entity F port map(lamdaA => P(9)(125),lamdaB => P(9)(127),lamdaOut => P(8)(125));
U_G9126: entity G port map(lamdaA => P(9)(124),lamdaB => P(9)(126),s => s(9)(62),lamdaOut => P(8)(126));
U_G9127: entity G port map(lamdaA => P(9)(125),lamdaB => P(9)(127),s => s(9)(63),lamdaOut => P(8)(127));
U_F9128: entity F port map(lamdaA => P(9)(128),lamdaB => P(9)(130),lamdaOut => P(8)(128));
U_F9129: entity F port map(lamdaA => P(9)(129),lamdaB => P(9)(131),lamdaOut => P(8)(129));
U_G9130: entity G port map(lamdaA => P(9)(128),lamdaB => P(9)(130),s => s(9)(64),lamdaOut => P(8)(130));
U_G9131: entity G port map(lamdaA => P(9)(129),lamdaB => P(9)(131),s => s(9)(65),lamdaOut => P(8)(131));
U_F9132: entity F port map(lamdaA => P(9)(132),lamdaB => P(9)(134),lamdaOut => P(8)(132));
U_F9133: entity F port map(lamdaA => P(9)(133),lamdaB => P(9)(135),lamdaOut => P(8)(133));
U_G9134: entity G port map(lamdaA => P(9)(132),lamdaB => P(9)(134),s => s(9)(66),lamdaOut => P(8)(134));
U_G9135: entity G port map(lamdaA => P(9)(133),lamdaB => P(9)(135),s => s(9)(67),lamdaOut => P(8)(135));
U_F9136: entity F port map(lamdaA => P(9)(136),lamdaB => P(9)(138),lamdaOut => P(8)(136));
U_F9137: entity F port map(lamdaA => P(9)(137),lamdaB => P(9)(139),lamdaOut => P(8)(137));
U_G9138: entity G port map(lamdaA => P(9)(136),lamdaB => P(9)(138),s => s(9)(68),lamdaOut => P(8)(138));
U_G9139: entity G port map(lamdaA => P(9)(137),lamdaB => P(9)(139),s => s(9)(69),lamdaOut => P(8)(139));
U_F9140: entity F port map(lamdaA => P(9)(140),lamdaB => P(9)(142),lamdaOut => P(8)(140));
U_F9141: entity F port map(lamdaA => P(9)(141),lamdaB => P(9)(143),lamdaOut => P(8)(141));
U_G9142: entity G port map(lamdaA => P(9)(140),lamdaB => P(9)(142),s => s(9)(70),lamdaOut => P(8)(142));
U_G9143: entity G port map(lamdaA => P(9)(141),lamdaB => P(9)(143),s => s(9)(71),lamdaOut => P(8)(143));
U_F9144: entity F port map(lamdaA => P(9)(144),lamdaB => P(9)(146),lamdaOut => P(8)(144));
U_F9145: entity F port map(lamdaA => P(9)(145),lamdaB => P(9)(147),lamdaOut => P(8)(145));
U_G9146: entity G port map(lamdaA => P(9)(144),lamdaB => P(9)(146),s => s(9)(72),lamdaOut => P(8)(146));
U_G9147: entity G port map(lamdaA => P(9)(145),lamdaB => P(9)(147),s => s(9)(73),lamdaOut => P(8)(147));
U_F9148: entity F port map(lamdaA => P(9)(148),lamdaB => P(9)(150),lamdaOut => P(8)(148));
U_F9149: entity F port map(lamdaA => P(9)(149),lamdaB => P(9)(151),lamdaOut => P(8)(149));
U_G9150: entity G port map(lamdaA => P(9)(148),lamdaB => P(9)(150),s => s(9)(74),lamdaOut => P(8)(150));
U_G9151: entity G port map(lamdaA => P(9)(149),lamdaB => P(9)(151),s => s(9)(75),lamdaOut => P(8)(151));
U_F9152: entity F port map(lamdaA => P(9)(152),lamdaB => P(9)(154),lamdaOut => P(8)(152));
U_F9153: entity F port map(lamdaA => P(9)(153),lamdaB => P(9)(155),lamdaOut => P(8)(153));
U_G9154: entity G port map(lamdaA => P(9)(152),lamdaB => P(9)(154),s => s(9)(76),lamdaOut => P(8)(154));
U_G9155: entity G port map(lamdaA => P(9)(153),lamdaB => P(9)(155),s => s(9)(77),lamdaOut => P(8)(155));
U_F9156: entity F port map(lamdaA => P(9)(156),lamdaB => P(9)(158),lamdaOut => P(8)(156));
U_F9157: entity F port map(lamdaA => P(9)(157),lamdaB => P(9)(159),lamdaOut => P(8)(157));
U_G9158: entity G port map(lamdaA => P(9)(156),lamdaB => P(9)(158),s => s(9)(78),lamdaOut => P(8)(158));
U_G9159: entity G port map(lamdaA => P(9)(157),lamdaB => P(9)(159),s => s(9)(79),lamdaOut => P(8)(159));
U_F9160: entity F port map(lamdaA => P(9)(160),lamdaB => P(9)(162),lamdaOut => P(8)(160));
U_F9161: entity F port map(lamdaA => P(9)(161),lamdaB => P(9)(163),lamdaOut => P(8)(161));
U_G9162: entity G port map(lamdaA => P(9)(160),lamdaB => P(9)(162),s => s(9)(80),lamdaOut => P(8)(162));
U_G9163: entity G port map(lamdaA => P(9)(161),lamdaB => P(9)(163),s => s(9)(81),lamdaOut => P(8)(163));
U_F9164: entity F port map(lamdaA => P(9)(164),lamdaB => P(9)(166),lamdaOut => P(8)(164));
U_F9165: entity F port map(lamdaA => P(9)(165),lamdaB => P(9)(167),lamdaOut => P(8)(165));
U_G9166: entity G port map(lamdaA => P(9)(164),lamdaB => P(9)(166),s => s(9)(82),lamdaOut => P(8)(166));
U_G9167: entity G port map(lamdaA => P(9)(165),lamdaB => P(9)(167),s => s(9)(83),lamdaOut => P(8)(167));
U_F9168: entity F port map(lamdaA => P(9)(168),lamdaB => P(9)(170),lamdaOut => P(8)(168));
U_F9169: entity F port map(lamdaA => P(9)(169),lamdaB => P(9)(171),lamdaOut => P(8)(169));
U_G9170: entity G port map(lamdaA => P(9)(168),lamdaB => P(9)(170),s => s(9)(84),lamdaOut => P(8)(170));
U_G9171: entity G port map(lamdaA => P(9)(169),lamdaB => P(9)(171),s => s(9)(85),lamdaOut => P(8)(171));
U_F9172: entity F port map(lamdaA => P(9)(172),lamdaB => P(9)(174),lamdaOut => P(8)(172));
U_F9173: entity F port map(lamdaA => P(9)(173),lamdaB => P(9)(175),lamdaOut => P(8)(173));
U_G9174: entity G port map(lamdaA => P(9)(172),lamdaB => P(9)(174),s => s(9)(86),lamdaOut => P(8)(174));
U_G9175: entity G port map(lamdaA => P(9)(173),lamdaB => P(9)(175),s => s(9)(87),lamdaOut => P(8)(175));
U_F9176: entity F port map(lamdaA => P(9)(176),lamdaB => P(9)(178),lamdaOut => P(8)(176));
U_F9177: entity F port map(lamdaA => P(9)(177),lamdaB => P(9)(179),lamdaOut => P(8)(177));
U_G9178: entity G port map(lamdaA => P(9)(176),lamdaB => P(9)(178),s => s(9)(88),lamdaOut => P(8)(178));
U_G9179: entity G port map(lamdaA => P(9)(177),lamdaB => P(9)(179),s => s(9)(89),lamdaOut => P(8)(179));
U_F9180: entity F port map(lamdaA => P(9)(180),lamdaB => P(9)(182),lamdaOut => P(8)(180));
U_F9181: entity F port map(lamdaA => P(9)(181),lamdaB => P(9)(183),lamdaOut => P(8)(181));
U_G9182: entity G port map(lamdaA => P(9)(180),lamdaB => P(9)(182),s => s(9)(90),lamdaOut => P(8)(182));
U_G9183: entity G port map(lamdaA => P(9)(181),lamdaB => P(9)(183),s => s(9)(91),lamdaOut => P(8)(183));
U_F9184: entity F port map(lamdaA => P(9)(184),lamdaB => P(9)(186),lamdaOut => P(8)(184));
U_F9185: entity F port map(lamdaA => P(9)(185),lamdaB => P(9)(187),lamdaOut => P(8)(185));
U_G9186: entity G port map(lamdaA => P(9)(184),lamdaB => P(9)(186),s => s(9)(92),lamdaOut => P(8)(186));
U_G9187: entity G port map(lamdaA => P(9)(185),lamdaB => P(9)(187),s => s(9)(93),lamdaOut => P(8)(187));
U_F9188: entity F port map(lamdaA => P(9)(188),lamdaB => P(9)(190),lamdaOut => P(8)(188));
U_F9189: entity F port map(lamdaA => P(9)(189),lamdaB => P(9)(191),lamdaOut => P(8)(189));
U_G9190: entity G port map(lamdaA => P(9)(188),lamdaB => P(9)(190),s => s(9)(94),lamdaOut => P(8)(190));
U_G9191: entity G port map(lamdaA => P(9)(189),lamdaB => P(9)(191),s => s(9)(95),lamdaOut => P(8)(191));
U_F9192: entity F port map(lamdaA => P(9)(192),lamdaB => P(9)(194),lamdaOut => P(8)(192));
U_F9193: entity F port map(lamdaA => P(9)(193),lamdaB => P(9)(195),lamdaOut => P(8)(193));
U_G9194: entity G port map(lamdaA => P(9)(192),lamdaB => P(9)(194),s => s(9)(96),lamdaOut => P(8)(194));
U_G9195: entity G port map(lamdaA => P(9)(193),lamdaB => P(9)(195),s => s(9)(97),lamdaOut => P(8)(195));
U_F9196: entity F port map(lamdaA => P(9)(196),lamdaB => P(9)(198),lamdaOut => P(8)(196));
U_F9197: entity F port map(lamdaA => P(9)(197),lamdaB => P(9)(199),lamdaOut => P(8)(197));
U_G9198: entity G port map(lamdaA => P(9)(196),lamdaB => P(9)(198),s => s(9)(98),lamdaOut => P(8)(198));
U_G9199: entity G port map(lamdaA => P(9)(197),lamdaB => P(9)(199),s => s(9)(99),lamdaOut => P(8)(199));
U_F9200: entity F port map(lamdaA => P(9)(200),lamdaB => P(9)(202),lamdaOut => P(8)(200));
U_F9201: entity F port map(lamdaA => P(9)(201),lamdaB => P(9)(203),lamdaOut => P(8)(201));
U_G9202: entity G port map(lamdaA => P(9)(200),lamdaB => P(9)(202),s => s(9)(100),lamdaOut => P(8)(202));
U_G9203: entity G port map(lamdaA => P(9)(201),lamdaB => P(9)(203),s => s(9)(101),lamdaOut => P(8)(203));
U_F9204: entity F port map(lamdaA => P(9)(204),lamdaB => P(9)(206),lamdaOut => P(8)(204));
U_F9205: entity F port map(lamdaA => P(9)(205),lamdaB => P(9)(207),lamdaOut => P(8)(205));
U_G9206: entity G port map(lamdaA => P(9)(204),lamdaB => P(9)(206),s => s(9)(102),lamdaOut => P(8)(206));
U_G9207: entity G port map(lamdaA => P(9)(205),lamdaB => P(9)(207),s => s(9)(103),lamdaOut => P(8)(207));
U_F9208: entity F port map(lamdaA => P(9)(208),lamdaB => P(9)(210),lamdaOut => P(8)(208));
U_F9209: entity F port map(lamdaA => P(9)(209),lamdaB => P(9)(211),lamdaOut => P(8)(209));
U_G9210: entity G port map(lamdaA => P(9)(208),lamdaB => P(9)(210),s => s(9)(104),lamdaOut => P(8)(210));
U_G9211: entity G port map(lamdaA => P(9)(209),lamdaB => P(9)(211),s => s(9)(105),lamdaOut => P(8)(211));
U_F9212: entity F port map(lamdaA => P(9)(212),lamdaB => P(9)(214),lamdaOut => P(8)(212));
U_F9213: entity F port map(lamdaA => P(9)(213),lamdaB => P(9)(215),lamdaOut => P(8)(213));
U_G9214: entity G port map(lamdaA => P(9)(212),lamdaB => P(9)(214),s => s(9)(106),lamdaOut => P(8)(214));
U_G9215: entity G port map(lamdaA => P(9)(213),lamdaB => P(9)(215),s => s(9)(107),lamdaOut => P(8)(215));
U_F9216: entity F port map(lamdaA => P(9)(216),lamdaB => P(9)(218),lamdaOut => P(8)(216));
U_F9217: entity F port map(lamdaA => P(9)(217),lamdaB => P(9)(219),lamdaOut => P(8)(217));
U_G9218: entity G port map(lamdaA => P(9)(216),lamdaB => P(9)(218),s => s(9)(108),lamdaOut => P(8)(218));
U_G9219: entity G port map(lamdaA => P(9)(217),lamdaB => P(9)(219),s => s(9)(109),lamdaOut => P(8)(219));
U_F9220: entity F port map(lamdaA => P(9)(220),lamdaB => P(9)(222),lamdaOut => P(8)(220));
U_F9221: entity F port map(lamdaA => P(9)(221),lamdaB => P(9)(223),lamdaOut => P(8)(221));
U_G9222: entity G port map(lamdaA => P(9)(220),lamdaB => P(9)(222),s => s(9)(110),lamdaOut => P(8)(222));
U_G9223: entity G port map(lamdaA => P(9)(221),lamdaB => P(9)(223),s => s(9)(111),lamdaOut => P(8)(223));
U_F9224: entity F port map(lamdaA => P(9)(224),lamdaB => P(9)(226),lamdaOut => P(8)(224));
U_F9225: entity F port map(lamdaA => P(9)(225),lamdaB => P(9)(227),lamdaOut => P(8)(225));
U_G9226: entity G port map(lamdaA => P(9)(224),lamdaB => P(9)(226),s => s(9)(112),lamdaOut => P(8)(226));
U_G9227: entity G port map(lamdaA => P(9)(225),lamdaB => P(9)(227),s => s(9)(113),lamdaOut => P(8)(227));
U_F9228: entity F port map(lamdaA => P(9)(228),lamdaB => P(9)(230),lamdaOut => P(8)(228));
U_F9229: entity F port map(lamdaA => P(9)(229),lamdaB => P(9)(231),lamdaOut => P(8)(229));
U_G9230: entity G port map(lamdaA => P(9)(228),lamdaB => P(9)(230),s => s(9)(114),lamdaOut => P(8)(230));
U_G9231: entity G port map(lamdaA => P(9)(229),lamdaB => P(9)(231),s => s(9)(115),lamdaOut => P(8)(231));
U_F9232: entity F port map(lamdaA => P(9)(232),lamdaB => P(9)(234),lamdaOut => P(8)(232));
U_F9233: entity F port map(lamdaA => P(9)(233),lamdaB => P(9)(235),lamdaOut => P(8)(233));
U_G9234: entity G port map(lamdaA => P(9)(232),lamdaB => P(9)(234),s => s(9)(116),lamdaOut => P(8)(234));
U_G9235: entity G port map(lamdaA => P(9)(233),lamdaB => P(9)(235),s => s(9)(117),lamdaOut => P(8)(235));
U_F9236: entity F port map(lamdaA => P(9)(236),lamdaB => P(9)(238),lamdaOut => P(8)(236));
U_F9237: entity F port map(lamdaA => P(9)(237),lamdaB => P(9)(239),lamdaOut => P(8)(237));
U_G9238: entity G port map(lamdaA => P(9)(236),lamdaB => P(9)(238),s => s(9)(118),lamdaOut => P(8)(238));
U_G9239: entity G port map(lamdaA => P(9)(237),lamdaB => P(9)(239),s => s(9)(119),lamdaOut => P(8)(239));
U_F9240: entity F port map(lamdaA => P(9)(240),lamdaB => P(9)(242),lamdaOut => P(8)(240));
U_F9241: entity F port map(lamdaA => P(9)(241),lamdaB => P(9)(243),lamdaOut => P(8)(241));
U_G9242: entity G port map(lamdaA => P(9)(240),lamdaB => P(9)(242),s => s(9)(120),lamdaOut => P(8)(242));
U_G9243: entity G port map(lamdaA => P(9)(241),lamdaB => P(9)(243),s => s(9)(121),lamdaOut => P(8)(243));
U_F9244: entity F port map(lamdaA => P(9)(244),lamdaB => P(9)(246),lamdaOut => P(8)(244));
U_F9245: entity F port map(lamdaA => P(9)(245),lamdaB => P(9)(247),lamdaOut => P(8)(245));
U_G9246: entity G port map(lamdaA => P(9)(244),lamdaB => P(9)(246),s => s(9)(122),lamdaOut => P(8)(246));
U_G9247: entity G port map(lamdaA => P(9)(245),lamdaB => P(9)(247),s => s(9)(123),lamdaOut => P(8)(247));
U_F9248: entity F port map(lamdaA => P(9)(248),lamdaB => P(9)(250),lamdaOut => P(8)(248));
U_F9249: entity F port map(lamdaA => P(9)(249),lamdaB => P(9)(251),lamdaOut => P(8)(249));
U_G9250: entity G port map(lamdaA => P(9)(248),lamdaB => P(9)(250),s => s(9)(124),lamdaOut => P(8)(250));
U_G9251: entity G port map(lamdaA => P(9)(249),lamdaB => P(9)(251),s => s(9)(125),lamdaOut => P(8)(251));
U_F9252: entity F port map(lamdaA => P(9)(252),lamdaB => P(9)(254),lamdaOut => P(8)(252));
U_F9253: entity F port map(lamdaA => P(9)(253),lamdaB => P(9)(255),lamdaOut => P(8)(253));
U_G9254: entity G port map(lamdaA => P(9)(252),lamdaB => P(9)(254),s => s(9)(126),lamdaOut => P(8)(254));
U_G9255: entity G port map(lamdaA => P(9)(253),lamdaB => P(9)(255),s => s(9)(127),lamdaOut => P(8)(255));
U_F9256: entity F port map(lamdaA => P(9)(256),lamdaB => P(9)(258),lamdaOut => P(8)(256));
U_F9257: entity F port map(lamdaA => P(9)(257),lamdaB => P(9)(259),lamdaOut => P(8)(257));
U_G9258: entity G port map(lamdaA => P(9)(256),lamdaB => P(9)(258),s => s(9)(128),lamdaOut => P(8)(258));
U_G9259: entity G port map(lamdaA => P(9)(257),lamdaB => P(9)(259),s => s(9)(129),lamdaOut => P(8)(259));
U_F9260: entity F port map(lamdaA => P(9)(260),lamdaB => P(9)(262),lamdaOut => P(8)(260));
U_F9261: entity F port map(lamdaA => P(9)(261),lamdaB => P(9)(263),lamdaOut => P(8)(261));
U_G9262: entity G port map(lamdaA => P(9)(260),lamdaB => P(9)(262),s => s(9)(130),lamdaOut => P(8)(262));
U_G9263: entity G port map(lamdaA => P(9)(261),lamdaB => P(9)(263),s => s(9)(131),lamdaOut => P(8)(263));
U_F9264: entity F port map(lamdaA => P(9)(264),lamdaB => P(9)(266),lamdaOut => P(8)(264));
U_F9265: entity F port map(lamdaA => P(9)(265),lamdaB => P(9)(267),lamdaOut => P(8)(265));
U_G9266: entity G port map(lamdaA => P(9)(264),lamdaB => P(9)(266),s => s(9)(132),lamdaOut => P(8)(266));
U_G9267: entity G port map(lamdaA => P(9)(265),lamdaB => P(9)(267),s => s(9)(133),lamdaOut => P(8)(267));
U_F9268: entity F port map(lamdaA => P(9)(268),lamdaB => P(9)(270),lamdaOut => P(8)(268));
U_F9269: entity F port map(lamdaA => P(9)(269),lamdaB => P(9)(271),lamdaOut => P(8)(269));
U_G9270: entity G port map(lamdaA => P(9)(268),lamdaB => P(9)(270),s => s(9)(134),lamdaOut => P(8)(270));
U_G9271: entity G port map(lamdaA => P(9)(269),lamdaB => P(9)(271),s => s(9)(135),lamdaOut => P(8)(271));
U_F9272: entity F port map(lamdaA => P(9)(272),lamdaB => P(9)(274),lamdaOut => P(8)(272));
U_F9273: entity F port map(lamdaA => P(9)(273),lamdaB => P(9)(275),lamdaOut => P(8)(273));
U_G9274: entity G port map(lamdaA => P(9)(272),lamdaB => P(9)(274),s => s(9)(136),lamdaOut => P(8)(274));
U_G9275: entity G port map(lamdaA => P(9)(273),lamdaB => P(9)(275),s => s(9)(137),lamdaOut => P(8)(275));
U_F9276: entity F port map(lamdaA => P(9)(276),lamdaB => P(9)(278),lamdaOut => P(8)(276));
U_F9277: entity F port map(lamdaA => P(9)(277),lamdaB => P(9)(279),lamdaOut => P(8)(277));
U_G9278: entity G port map(lamdaA => P(9)(276),lamdaB => P(9)(278),s => s(9)(138),lamdaOut => P(8)(278));
U_G9279: entity G port map(lamdaA => P(9)(277),lamdaB => P(9)(279),s => s(9)(139),lamdaOut => P(8)(279));
U_F9280: entity F port map(lamdaA => P(9)(280),lamdaB => P(9)(282),lamdaOut => P(8)(280));
U_F9281: entity F port map(lamdaA => P(9)(281),lamdaB => P(9)(283),lamdaOut => P(8)(281));
U_G9282: entity G port map(lamdaA => P(9)(280),lamdaB => P(9)(282),s => s(9)(140),lamdaOut => P(8)(282));
U_G9283: entity G port map(lamdaA => P(9)(281),lamdaB => P(9)(283),s => s(9)(141),lamdaOut => P(8)(283));
U_F9284: entity F port map(lamdaA => P(9)(284),lamdaB => P(9)(286),lamdaOut => P(8)(284));
U_F9285: entity F port map(lamdaA => P(9)(285),lamdaB => P(9)(287),lamdaOut => P(8)(285));
U_G9286: entity G port map(lamdaA => P(9)(284),lamdaB => P(9)(286),s => s(9)(142),lamdaOut => P(8)(286));
U_G9287: entity G port map(lamdaA => P(9)(285),lamdaB => P(9)(287),s => s(9)(143),lamdaOut => P(8)(287));
U_F9288: entity F port map(lamdaA => P(9)(288),lamdaB => P(9)(290),lamdaOut => P(8)(288));
U_F9289: entity F port map(lamdaA => P(9)(289),lamdaB => P(9)(291),lamdaOut => P(8)(289));
U_G9290: entity G port map(lamdaA => P(9)(288),lamdaB => P(9)(290),s => s(9)(144),lamdaOut => P(8)(290));
U_G9291: entity G port map(lamdaA => P(9)(289),lamdaB => P(9)(291),s => s(9)(145),lamdaOut => P(8)(291));
U_F9292: entity F port map(lamdaA => P(9)(292),lamdaB => P(9)(294),lamdaOut => P(8)(292));
U_F9293: entity F port map(lamdaA => P(9)(293),lamdaB => P(9)(295),lamdaOut => P(8)(293));
U_G9294: entity G port map(lamdaA => P(9)(292),lamdaB => P(9)(294),s => s(9)(146),lamdaOut => P(8)(294));
U_G9295: entity G port map(lamdaA => P(9)(293),lamdaB => P(9)(295),s => s(9)(147),lamdaOut => P(8)(295));
U_F9296: entity F port map(lamdaA => P(9)(296),lamdaB => P(9)(298),lamdaOut => P(8)(296));
U_F9297: entity F port map(lamdaA => P(9)(297),lamdaB => P(9)(299),lamdaOut => P(8)(297));
U_G9298: entity G port map(lamdaA => P(9)(296),lamdaB => P(9)(298),s => s(9)(148),lamdaOut => P(8)(298));
U_G9299: entity G port map(lamdaA => P(9)(297),lamdaB => P(9)(299),s => s(9)(149),lamdaOut => P(8)(299));
U_F9300: entity F port map(lamdaA => P(9)(300),lamdaB => P(9)(302),lamdaOut => P(8)(300));
U_F9301: entity F port map(lamdaA => P(9)(301),lamdaB => P(9)(303),lamdaOut => P(8)(301));
U_G9302: entity G port map(lamdaA => P(9)(300),lamdaB => P(9)(302),s => s(9)(150),lamdaOut => P(8)(302));
U_G9303: entity G port map(lamdaA => P(9)(301),lamdaB => P(9)(303),s => s(9)(151),lamdaOut => P(8)(303));
U_F9304: entity F port map(lamdaA => P(9)(304),lamdaB => P(9)(306),lamdaOut => P(8)(304));
U_F9305: entity F port map(lamdaA => P(9)(305),lamdaB => P(9)(307),lamdaOut => P(8)(305));
U_G9306: entity G port map(lamdaA => P(9)(304),lamdaB => P(9)(306),s => s(9)(152),lamdaOut => P(8)(306));
U_G9307: entity G port map(lamdaA => P(9)(305),lamdaB => P(9)(307),s => s(9)(153),lamdaOut => P(8)(307));
U_F9308: entity F port map(lamdaA => P(9)(308),lamdaB => P(9)(310),lamdaOut => P(8)(308));
U_F9309: entity F port map(lamdaA => P(9)(309),lamdaB => P(9)(311),lamdaOut => P(8)(309));
U_G9310: entity G port map(lamdaA => P(9)(308),lamdaB => P(9)(310),s => s(9)(154),lamdaOut => P(8)(310));
U_G9311: entity G port map(lamdaA => P(9)(309),lamdaB => P(9)(311),s => s(9)(155),lamdaOut => P(8)(311));
U_F9312: entity F port map(lamdaA => P(9)(312),lamdaB => P(9)(314),lamdaOut => P(8)(312));
U_F9313: entity F port map(lamdaA => P(9)(313),lamdaB => P(9)(315),lamdaOut => P(8)(313));
U_G9314: entity G port map(lamdaA => P(9)(312),lamdaB => P(9)(314),s => s(9)(156),lamdaOut => P(8)(314));
U_G9315: entity G port map(lamdaA => P(9)(313),lamdaB => P(9)(315),s => s(9)(157),lamdaOut => P(8)(315));
U_F9316: entity F port map(lamdaA => P(9)(316),lamdaB => P(9)(318),lamdaOut => P(8)(316));
U_F9317: entity F port map(lamdaA => P(9)(317),lamdaB => P(9)(319),lamdaOut => P(8)(317));
U_G9318: entity G port map(lamdaA => P(9)(316),lamdaB => P(9)(318),s => s(9)(158),lamdaOut => P(8)(318));
U_G9319: entity G port map(lamdaA => P(9)(317),lamdaB => P(9)(319),s => s(9)(159),lamdaOut => P(8)(319));
U_F9320: entity F port map(lamdaA => P(9)(320),lamdaB => P(9)(322),lamdaOut => P(8)(320));
U_F9321: entity F port map(lamdaA => P(9)(321),lamdaB => P(9)(323),lamdaOut => P(8)(321));
U_G9322: entity G port map(lamdaA => P(9)(320),lamdaB => P(9)(322),s => s(9)(160),lamdaOut => P(8)(322));
U_G9323: entity G port map(lamdaA => P(9)(321),lamdaB => P(9)(323),s => s(9)(161),lamdaOut => P(8)(323));
U_F9324: entity F port map(lamdaA => P(9)(324),lamdaB => P(9)(326),lamdaOut => P(8)(324));
U_F9325: entity F port map(lamdaA => P(9)(325),lamdaB => P(9)(327),lamdaOut => P(8)(325));
U_G9326: entity G port map(lamdaA => P(9)(324),lamdaB => P(9)(326),s => s(9)(162),lamdaOut => P(8)(326));
U_G9327: entity G port map(lamdaA => P(9)(325),lamdaB => P(9)(327),s => s(9)(163),lamdaOut => P(8)(327));
U_F9328: entity F port map(lamdaA => P(9)(328),lamdaB => P(9)(330),lamdaOut => P(8)(328));
U_F9329: entity F port map(lamdaA => P(9)(329),lamdaB => P(9)(331),lamdaOut => P(8)(329));
U_G9330: entity G port map(lamdaA => P(9)(328),lamdaB => P(9)(330),s => s(9)(164),lamdaOut => P(8)(330));
U_G9331: entity G port map(lamdaA => P(9)(329),lamdaB => P(9)(331),s => s(9)(165),lamdaOut => P(8)(331));
U_F9332: entity F port map(lamdaA => P(9)(332),lamdaB => P(9)(334),lamdaOut => P(8)(332));
U_F9333: entity F port map(lamdaA => P(9)(333),lamdaB => P(9)(335),lamdaOut => P(8)(333));
U_G9334: entity G port map(lamdaA => P(9)(332),lamdaB => P(9)(334),s => s(9)(166),lamdaOut => P(8)(334));
U_G9335: entity G port map(lamdaA => P(9)(333),lamdaB => P(9)(335),s => s(9)(167),lamdaOut => P(8)(335));
U_F9336: entity F port map(lamdaA => P(9)(336),lamdaB => P(9)(338),lamdaOut => P(8)(336));
U_F9337: entity F port map(lamdaA => P(9)(337),lamdaB => P(9)(339),lamdaOut => P(8)(337));
U_G9338: entity G port map(lamdaA => P(9)(336),lamdaB => P(9)(338),s => s(9)(168),lamdaOut => P(8)(338));
U_G9339: entity G port map(lamdaA => P(9)(337),lamdaB => P(9)(339),s => s(9)(169),lamdaOut => P(8)(339));
U_F9340: entity F port map(lamdaA => P(9)(340),lamdaB => P(9)(342),lamdaOut => P(8)(340));
U_F9341: entity F port map(lamdaA => P(9)(341),lamdaB => P(9)(343),lamdaOut => P(8)(341));
U_G9342: entity G port map(lamdaA => P(9)(340),lamdaB => P(9)(342),s => s(9)(170),lamdaOut => P(8)(342));
U_G9343: entity G port map(lamdaA => P(9)(341),lamdaB => P(9)(343),s => s(9)(171),lamdaOut => P(8)(343));
U_F9344: entity F port map(lamdaA => P(9)(344),lamdaB => P(9)(346),lamdaOut => P(8)(344));
U_F9345: entity F port map(lamdaA => P(9)(345),lamdaB => P(9)(347),lamdaOut => P(8)(345));
U_G9346: entity G port map(lamdaA => P(9)(344),lamdaB => P(9)(346),s => s(9)(172),lamdaOut => P(8)(346));
U_G9347: entity G port map(lamdaA => P(9)(345),lamdaB => P(9)(347),s => s(9)(173),lamdaOut => P(8)(347));
U_F9348: entity F port map(lamdaA => P(9)(348),lamdaB => P(9)(350),lamdaOut => P(8)(348));
U_F9349: entity F port map(lamdaA => P(9)(349),lamdaB => P(9)(351),lamdaOut => P(8)(349));
U_G9350: entity G port map(lamdaA => P(9)(348),lamdaB => P(9)(350),s => s(9)(174),lamdaOut => P(8)(350));
U_G9351: entity G port map(lamdaA => P(9)(349),lamdaB => P(9)(351),s => s(9)(175),lamdaOut => P(8)(351));
U_F9352: entity F port map(lamdaA => P(9)(352),lamdaB => P(9)(354),lamdaOut => P(8)(352));
U_F9353: entity F port map(lamdaA => P(9)(353),lamdaB => P(9)(355),lamdaOut => P(8)(353));
U_G9354: entity G port map(lamdaA => P(9)(352),lamdaB => P(9)(354),s => s(9)(176),lamdaOut => P(8)(354));
U_G9355: entity G port map(lamdaA => P(9)(353),lamdaB => P(9)(355),s => s(9)(177),lamdaOut => P(8)(355));
U_F9356: entity F port map(lamdaA => P(9)(356),lamdaB => P(9)(358),lamdaOut => P(8)(356));
U_F9357: entity F port map(lamdaA => P(9)(357),lamdaB => P(9)(359),lamdaOut => P(8)(357));
U_G9358: entity G port map(lamdaA => P(9)(356),lamdaB => P(9)(358),s => s(9)(178),lamdaOut => P(8)(358));
U_G9359: entity G port map(lamdaA => P(9)(357),lamdaB => P(9)(359),s => s(9)(179),lamdaOut => P(8)(359));
U_F9360: entity F port map(lamdaA => P(9)(360),lamdaB => P(9)(362),lamdaOut => P(8)(360));
U_F9361: entity F port map(lamdaA => P(9)(361),lamdaB => P(9)(363),lamdaOut => P(8)(361));
U_G9362: entity G port map(lamdaA => P(9)(360),lamdaB => P(9)(362),s => s(9)(180),lamdaOut => P(8)(362));
U_G9363: entity G port map(lamdaA => P(9)(361),lamdaB => P(9)(363),s => s(9)(181),lamdaOut => P(8)(363));
U_F9364: entity F port map(lamdaA => P(9)(364),lamdaB => P(9)(366),lamdaOut => P(8)(364));
U_F9365: entity F port map(lamdaA => P(9)(365),lamdaB => P(9)(367),lamdaOut => P(8)(365));
U_G9366: entity G port map(lamdaA => P(9)(364),lamdaB => P(9)(366),s => s(9)(182),lamdaOut => P(8)(366));
U_G9367: entity G port map(lamdaA => P(9)(365),lamdaB => P(9)(367),s => s(9)(183),lamdaOut => P(8)(367));
U_F9368: entity F port map(lamdaA => P(9)(368),lamdaB => P(9)(370),lamdaOut => P(8)(368));
U_F9369: entity F port map(lamdaA => P(9)(369),lamdaB => P(9)(371),lamdaOut => P(8)(369));
U_G9370: entity G port map(lamdaA => P(9)(368),lamdaB => P(9)(370),s => s(9)(184),lamdaOut => P(8)(370));
U_G9371: entity G port map(lamdaA => P(9)(369),lamdaB => P(9)(371),s => s(9)(185),lamdaOut => P(8)(371));
U_F9372: entity F port map(lamdaA => P(9)(372),lamdaB => P(9)(374),lamdaOut => P(8)(372));
U_F9373: entity F port map(lamdaA => P(9)(373),lamdaB => P(9)(375),lamdaOut => P(8)(373));
U_G9374: entity G port map(lamdaA => P(9)(372),lamdaB => P(9)(374),s => s(9)(186),lamdaOut => P(8)(374));
U_G9375: entity G port map(lamdaA => P(9)(373),lamdaB => P(9)(375),s => s(9)(187),lamdaOut => P(8)(375));
U_F9376: entity F port map(lamdaA => P(9)(376),lamdaB => P(9)(378),lamdaOut => P(8)(376));
U_F9377: entity F port map(lamdaA => P(9)(377),lamdaB => P(9)(379),lamdaOut => P(8)(377));
U_G9378: entity G port map(lamdaA => P(9)(376),lamdaB => P(9)(378),s => s(9)(188),lamdaOut => P(8)(378));
U_G9379: entity G port map(lamdaA => P(9)(377),lamdaB => P(9)(379),s => s(9)(189),lamdaOut => P(8)(379));
U_F9380: entity F port map(lamdaA => P(9)(380),lamdaB => P(9)(382),lamdaOut => P(8)(380));
U_F9381: entity F port map(lamdaA => P(9)(381),lamdaB => P(9)(383),lamdaOut => P(8)(381));
U_G9382: entity G port map(lamdaA => P(9)(380),lamdaB => P(9)(382),s => s(9)(190),lamdaOut => P(8)(382));
U_G9383: entity G port map(lamdaA => P(9)(381),lamdaB => P(9)(383),s => s(9)(191),lamdaOut => P(8)(383));
U_F9384: entity F port map(lamdaA => P(9)(384),lamdaB => P(9)(386),lamdaOut => P(8)(384));
U_F9385: entity F port map(lamdaA => P(9)(385),lamdaB => P(9)(387),lamdaOut => P(8)(385));
U_G9386: entity G port map(lamdaA => P(9)(384),lamdaB => P(9)(386),s => s(9)(192),lamdaOut => P(8)(386));
U_G9387: entity G port map(lamdaA => P(9)(385),lamdaB => P(9)(387),s => s(9)(193),lamdaOut => P(8)(387));
U_F9388: entity F port map(lamdaA => P(9)(388),lamdaB => P(9)(390),lamdaOut => P(8)(388));
U_F9389: entity F port map(lamdaA => P(9)(389),lamdaB => P(9)(391),lamdaOut => P(8)(389));
U_G9390: entity G port map(lamdaA => P(9)(388),lamdaB => P(9)(390),s => s(9)(194),lamdaOut => P(8)(390));
U_G9391: entity G port map(lamdaA => P(9)(389),lamdaB => P(9)(391),s => s(9)(195),lamdaOut => P(8)(391));
U_F9392: entity F port map(lamdaA => P(9)(392),lamdaB => P(9)(394),lamdaOut => P(8)(392));
U_F9393: entity F port map(lamdaA => P(9)(393),lamdaB => P(9)(395),lamdaOut => P(8)(393));
U_G9394: entity G port map(lamdaA => P(9)(392),lamdaB => P(9)(394),s => s(9)(196),lamdaOut => P(8)(394));
U_G9395: entity G port map(lamdaA => P(9)(393),lamdaB => P(9)(395),s => s(9)(197),lamdaOut => P(8)(395));
U_F9396: entity F port map(lamdaA => P(9)(396),lamdaB => P(9)(398),lamdaOut => P(8)(396));
U_F9397: entity F port map(lamdaA => P(9)(397),lamdaB => P(9)(399),lamdaOut => P(8)(397));
U_G9398: entity G port map(lamdaA => P(9)(396),lamdaB => P(9)(398),s => s(9)(198),lamdaOut => P(8)(398));
U_G9399: entity G port map(lamdaA => P(9)(397),lamdaB => P(9)(399),s => s(9)(199),lamdaOut => P(8)(399));
U_F9400: entity F port map(lamdaA => P(9)(400),lamdaB => P(9)(402),lamdaOut => P(8)(400));
U_F9401: entity F port map(lamdaA => P(9)(401),lamdaB => P(9)(403),lamdaOut => P(8)(401));
U_G9402: entity G port map(lamdaA => P(9)(400),lamdaB => P(9)(402),s => s(9)(200),lamdaOut => P(8)(402));
U_G9403: entity G port map(lamdaA => P(9)(401),lamdaB => P(9)(403),s => s(9)(201),lamdaOut => P(8)(403));
U_F9404: entity F port map(lamdaA => P(9)(404),lamdaB => P(9)(406),lamdaOut => P(8)(404));
U_F9405: entity F port map(lamdaA => P(9)(405),lamdaB => P(9)(407),lamdaOut => P(8)(405));
U_G9406: entity G port map(lamdaA => P(9)(404),lamdaB => P(9)(406),s => s(9)(202),lamdaOut => P(8)(406));
U_G9407: entity G port map(lamdaA => P(9)(405),lamdaB => P(9)(407),s => s(9)(203),lamdaOut => P(8)(407));
U_F9408: entity F port map(lamdaA => P(9)(408),lamdaB => P(9)(410),lamdaOut => P(8)(408));
U_F9409: entity F port map(lamdaA => P(9)(409),lamdaB => P(9)(411),lamdaOut => P(8)(409));
U_G9410: entity G port map(lamdaA => P(9)(408),lamdaB => P(9)(410),s => s(9)(204),lamdaOut => P(8)(410));
U_G9411: entity G port map(lamdaA => P(9)(409),lamdaB => P(9)(411),s => s(9)(205),lamdaOut => P(8)(411));
U_F9412: entity F port map(lamdaA => P(9)(412),lamdaB => P(9)(414),lamdaOut => P(8)(412));
U_F9413: entity F port map(lamdaA => P(9)(413),lamdaB => P(9)(415),lamdaOut => P(8)(413));
U_G9414: entity G port map(lamdaA => P(9)(412),lamdaB => P(9)(414),s => s(9)(206),lamdaOut => P(8)(414));
U_G9415: entity G port map(lamdaA => P(9)(413),lamdaB => P(9)(415),s => s(9)(207),lamdaOut => P(8)(415));
U_F9416: entity F port map(lamdaA => P(9)(416),lamdaB => P(9)(418),lamdaOut => P(8)(416));
U_F9417: entity F port map(lamdaA => P(9)(417),lamdaB => P(9)(419),lamdaOut => P(8)(417));
U_G9418: entity G port map(lamdaA => P(9)(416),lamdaB => P(9)(418),s => s(9)(208),lamdaOut => P(8)(418));
U_G9419: entity G port map(lamdaA => P(9)(417),lamdaB => P(9)(419),s => s(9)(209),lamdaOut => P(8)(419));
U_F9420: entity F port map(lamdaA => P(9)(420),lamdaB => P(9)(422),lamdaOut => P(8)(420));
U_F9421: entity F port map(lamdaA => P(9)(421),lamdaB => P(9)(423),lamdaOut => P(8)(421));
U_G9422: entity G port map(lamdaA => P(9)(420),lamdaB => P(9)(422),s => s(9)(210),lamdaOut => P(8)(422));
U_G9423: entity G port map(lamdaA => P(9)(421),lamdaB => P(9)(423),s => s(9)(211),lamdaOut => P(8)(423));
U_F9424: entity F port map(lamdaA => P(9)(424),lamdaB => P(9)(426),lamdaOut => P(8)(424));
U_F9425: entity F port map(lamdaA => P(9)(425),lamdaB => P(9)(427),lamdaOut => P(8)(425));
U_G9426: entity G port map(lamdaA => P(9)(424),lamdaB => P(9)(426),s => s(9)(212),lamdaOut => P(8)(426));
U_G9427: entity G port map(lamdaA => P(9)(425),lamdaB => P(9)(427),s => s(9)(213),lamdaOut => P(8)(427));
U_F9428: entity F port map(lamdaA => P(9)(428),lamdaB => P(9)(430),lamdaOut => P(8)(428));
U_F9429: entity F port map(lamdaA => P(9)(429),lamdaB => P(9)(431),lamdaOut => P(8)(429));
U_G9430: entity G port map(lamdaA => P(9)(428),lamdaB => P(9)(430),s => s(9)(214),lamdaOut => P(8)(430));
U_G9431: entity G port map(lamdaA => P(9)(429),lamdaB => P(9)(431),s => s(9)(215),lamdaOut => P(8)(431));
U_F9432: entity F port map(lamdaA => P(9)(432),lamdaB => P(9)(434),lamdaOut => P(8)(432));
U_F9433: entity F port map(lamdaA => P(9)(433),lamdaB => P(9)(435),lamdaOut => P(8)(433));
U_G9434: entity G port map(lamdaA => P(9)(432),lamdaB => P(9)(434),s => s(9)(216),lamdaOut => P(8)(434));
U_G9435: entity G port map(lamdaA => P(9)(433),lamdaB => P(9)(435),s => s(9)(217),lamdaOut => P(8)(435));
U_F9436: entity F port map(lamdaA => P(9)(436),lamdaB => P(9)(438),lamdaOut => P(8)(436));
U_F9437: entity F port map(lamdaA => P(9)(437),lamdaB => P(9)(439),lamdaOut => P(8)(437));
U_G9438: entity G port map(lamdaA => P(9)(436),lamdaB => P(9)(438),s => s(9)(218),lamdaOut => P(8)(438));
U_G9439: entity G port map(lamdaA => P(9)(437),lamdaB => P(9)(439),s => s(9)(219),lamdaOut => P(8)(439));
U_F9440: entity F port map(lamdaA => P(9)(440),lamdaB => P(9)(442),lamdaOut => P(8)(440));
U_F9441: entity F port map(lamdaA => P(9)(441),lamdaB => P(9)(443),lamdaOut => P(8)(441));
U_G9442: entity G port map(lamdaA => P(9)(440),lamdaB => P(9)(442),s => s(9)(220),lamdaOut => P(8)(442));
U_G9443: entity G port map(lamdaA => P(9)(441),lamdaB => P(9)(443),s => s(9)(221),lamdaOut => P(8)(443));
U_F9444: entity F port map(lamdaA => P(9)(444),lamdaB => P(9)(446),lamdaOut => P(8)(444));
U_F9445: entity F port map(lamdaA => P(9)(445),lamdaB => P(9)(447),lamdaOut => P(8)(445));
U_G9446: entity G port map(lamdaA => P(9)(444),lamdaB => P(9)(446),s => s(9)(222),lamdaOut => P(8)(446));
U_G9447: entity G port map(lamdaA => P(9)(445),lamdaB => P(9)(447),s => s(9)(223),lamdaOut => P(8)(447));
U_F9448: entity F port map(lamdaA => P(9)(448),lamdaB => P(9)(450),lamdaOut => P(8)(448));
U_F9449: entity F port map(lamdaA => P(9)(449),lamdaB => P(9)(451),lamdaOut => P(8)(449));
U_G9450: entity G port map(lamdaA => P(9)(448),lamdaB => P(9)(450),s => s(9)(224),lamdaOut => P(8)(450));
U_G9451: entity G port map(lamdaA => P(9)(449),lamdaB => P(9)(451),s => s(9)(225),lamdaOut => P(8)(451));
U_F9452: entity F port map(lamdaA => P(9)(452),lamdaB => P(9)(454),lamdaOut => P(8)(452));
U_F9453: entity F port map(lamdaA => P(9)(453),lamdaB => P(9)(455),lamdaOut => P(8)(453));
U_G9454: entity G port map(lamdaA => P(9)(452),lamdaB => P(9)(454),s => s(9)(226),lamdaOut => P(8)(454));
U_G9455: entity G port map(lamdaA => P(9)(453),lamdaB => P(9)(455),s => s(9)(227),lamdaOut => P(8)(455));
U_F9456: entity F port map(lamdaA => P(9)(456),lamdaB => P(9)(458),lamdaOut => P(8)(456));
U_F9457: entity F port map(lamdaA => P(9)(457),lamdaB => P(9)(459),lamdaOut => P(8)(457));
U_G9458: entity G port map(lamdaA => P(9)(456),lamdaB => P(9)(458),s => s(9)(228),lamdaOut => P(8)(458));
U_G9459: entity G port map(lamdaA => P(9)(457),lamdaB => P(9)(459),s => s(9)(229),lamdaOut => P(8)(459));
U_F9460: entity F port map(lamdaA => P(9)(460),lamdaB => P(9)(462),lamdaOut => P(8)(460));
U_F9461: entity F port map(lamdaA => P(9)(461),lamdaB => P(9)(463),lamdaOut => P(8)(461));
U_G9462: entity G port map(lamdaA => P(9)(460),lamdaB => P(9)(462),s => s(9)(230),lamdaOut => P(8)(462));
U_G9463: entity G port map(lamdaA => P(9)(461),lamdaB => P(9)(463),s => s(9)(231),lamdaOut => P(8)(463));
U_F9464: entity F port map(lamdaA => P(9)(464),lamdaB => P(9)(466),lamdaOut => P(8)(464));
U_F9465: entity F port map(lamdaA => P(9)(465),lamdaB => P(9)(467),lamdaOut => P(8)(465));
U_G9466: entity G port map(lamdaA => P(9)(464),lamdaB => P(9)(466),s => s(9)(232),lamdaOut => P(8)(466));
U_G9467: entity G port map(lamdaA => P(9)(465),lamdaB => P(9)(467),s => s(9)(233),lamdaOut => P(8)(467));
U_F9468: entity F port map(lamdaA => P(9)(468),lamdaB => P(9)(470),lamdaOut => P(8)(468));
U_F9469: entity F port map(lamdaA => P(9)(469),lamdaB => P(9)(471),lamdaOut => P(8)(469));
U_G9470: entity G port map(lamdaA => P(9)(468),lamdaB => P(9)(470),s => s(9)(234),lamdaOut => P(8)(470));
U_G9471: entity G port map(lamdaA => P(9)(469),lamdaB => P(9)(471),s => s(9)(235),lamdaOut => P(8)(471));
U_F9472: entity F port map(lamdaA => P(9)(472),lamdaB => P(9)(474),lamdaOut => P(8)(472));
U_F9473: entity F port map(lamdaA => P(9)(473),lamdaB => P(9)(475),lamdaOut => P(8)(473));
U_G9474: entity G port map(lamdaA => P(9)(472),lamdaB => P(9)(474),s => s(9)(236),lamdaOut => P(8)(474));
U_G9475: entity G port map(lamdaA => P(9)(473),lamdaB => P(9)(475),s => s(9)(237),lamdaOut => P(8)(475));
U_F9476: entity F port map(lamdaA => P(9)(476),lamdaB => P(9)(478),lamdaOut => P(8)(476));
U_F9477: entity F port map(lamdaA => P(9)(477),lamdaB => P(9)(479),lamdaOut => P(8)(477));
U_G9478: entity G port map(lamdaA => P(9)(476),lamdaB => P(9)(478),s => s(9)(238),lamdaOut => P(8)(478));
U_G9479: entity G port map(lamdaA => P(9)(477),lamdaB => P(9)(479),s => s(9)(239),lamdaOut => P(8)(479));
U_F9480: entity F port map(lamdaA => P(9)(480),lamdaB => P(9)(482),lamdaOut => P(8)(480));
U_F9481: entity F port map(lamdaA => P(9)(481),lamdaB => P(9)(483),lamdaOut => P(8)(481));
U_G9482: entity G port map(lamdaA => P(9)(480),lamdaB => P(9)(482),s => s(9)(240),lamdaOut => P(8)(482));
U_G9483: entity G port map(lamdaA => P(9)(481),lamdaB => P(9)(483),s => s(9)(241),lamdaOut => P(8)(483));
U_F9484: entity F port map(lamdaA => P(9)(484),lamdaB => P(9)(486),lamdaOut => P(8)(484));
U_F9485: entity F port map(lamdaA => P(9)(485),lamdaB => P(9)(487),lamdaOut => P(8)(485));
U_G9486: entity G port map(lamdaA => P(9)(484),lamdaB => P(9)(486),s => s(9)(242),lamdaOut => P(8)(486));
U_G9487: entity G port map(lamdaA => P(9)(485),lamdaB => P(9)(487),s => s(9)(243),lamdaOut => P(8)(487));
U_F9488: entity F port map(lamdaA => P(9)(488),lamdaB => P(9)(490),lamdaOut => P(8)(488));
U_F9489: entity F port map(lamdaA => P(9)(489),lamdaB => P(9)(491),lamdaOut => P(8)(489));
U_G9490: entity G port map(lamdaA => P(9)(488),lamdaB => P(9)(490),s => s(9)(244),lamdaOut => P(8)(490));
U_G9491: entity G port map(lamdaA => P(9)(489),lamdaB => P(9)(491),s => s(9)(245),lamdaOut => P(8)(491));
U_F9492: entity F port map(lamdaA => P(9)(492),lamdaB => P(9)(494),lamdaOut => P(8)(492));
U_F9493: entity F port map(lamdaA => P(9)(493),lamdaB => P(9)(495),lamdaOut => P(8)(493));
U_G9494: entity G port map(lamdaA => P(9)(492),lamdaB => P(9)(494),s => s(9)(246),lamdaOut => P(8)(494));
U_G9495: entity G port map(lamdaA => P(9)(493),lamdaB => P(9)(495),s => s(9)(247),lamdaOut => P(8)(495));
U_F9496: entity F port map(lamdaA => P(9)(496),lamdaB => P(9)(498),lamdaOut => P(8)(496));
U_F9497: entity F port map(lamdaA => P(9)(497),lamdaB => P(9)(499),lamdaOut => P(8)(497));
U_G9498: entity G port map(lamdaA => P(9)(496),lamdaB => P(9)(498),s => s(9)(248),lamdaOut => P(8)(498));
U_G9499: entity G port map(lamdaA => P(9)(497),lamdaB => P(9)(499),s => s(9)(249),lamdaOut => P(8)(499));
U_F9500: entity F port map(lamdaA => P(9)(500),lamdaB => P(9)(502),lamdaOut => P(8)(500));
U_F9501: entity F port map(lamdaA => P(9)(501),lamdaB => P(9)(503),lamdaOut => P(8)(501));
U_G9502: entity G port map(lamdaA => P(9)(500),lamdaB => P(9)(502),s => s(9)(250),lamdaOut => P(8)(502));
U_G9503: entity G port map(lamdaA => P(9)(501),lamdaB => P(9)(503),s => s(9)(251),lamdaOut => P(8)(503));
U_F9504: entity F port map(lamdaA => P(9)(504),lamdaB => P(9)(506),lamdaOut => P(8)(504));
U_F9505: entity F port map(lamdaA => P(9)(505),lamdaB => P(9)(507),lamdaOut => P(8)(505));
U_G9506: entity G port map(lamdaA => P(9)(504),lamdaB => P(9)(506),s => s(9)(252),lamdaOut => P(8)(506));
U_G9507: entity G port map(lamdaA => P(9)(505),lamdaB => P(9)(507),s => s(9)(253),lamdaOut => P(8)(507));
U_F9508: entity F port map(lamdaA => P(9)(508),lamdaB => P(9)(510),lamdaOut => P(8)(508));
U_F9509: entity F port map(lamdaA => P(9)(509),lamdaB => P(9)(511),lamdaOut => P(8)(509));
U_G9510: entity G port map(lamdaA => P(9)(508),lamdaB => P(9)(510),s => s(9)(254),lamdaOut => P(8)(510));
U_G9511: entity G port map(lamdaA => P(9)(509),lamdaB => P(9)(511),s => s(9)(255),lamdaOut => P(8)(511));
U_F9512: entity F port map(lamdaA => P(9)(512),lamdaB => P(9)(514),lamdaOut => P(8)(512));
U_F9513: entity F port map(lamdaA => P(9)(513),lamdaB => P(9)(515),lamdaOut => P(8)(513));
U_G9514: entity G port map(lamdaA => P(9)(512),lamdaB => P(9)(514),s => s(9)(256),lamdaOut => P(8)(514));
U_G9515: entity G port map(lamdaA => P(9)(513),lamdaB => P(9)(515),s => s(9)(257),lamdaOut => P(8)(515));
U_F9516: entity F port map(lamdaA => P(9)(516),lamdaB => P(9)(518),lamdaOut => P(8)(516));
U_F9517: entity F port map(lamdaA => P(9)(517),lamdaB => P(9)(519),lamdaOut => P(8)(517));
U_G9518: entity G port map(lamdaA => P(9)(516),lamdaB => P(9)(518),s => s(9)(258),lamdaOut => P(8)(518));
U_G9519: entity G port map(lamdaA => P(9)(517),lamdaB => P(9)(519),s => s(9)(259),lamdaOut => P(8)(519));
U_F9520: entity F port map(lamdaA => P(9)(520),lamdaB => P(9)(522),lamdaOut => P(8)(520));
U_F9521: entity F port map(lamdaA => P(9)(521),lamdaB => P(9)(523),lamdaOut => P(8)(521));
U_G9522: entity G port map(lamdaA => P(9)(520),lamdaB => P(9)(522),s => s(9)(260),lamdaOut => P(8)(522));
U_G9523: entity G port map(lamdaA => P(9)(521),lamdaB => P(9)(523),s => s(9)(261),lamdaOut => P(8)(523));
U_F9524: entity F port map(lamdaA => P(9)(524),lamdaB => P(9)(526),lamdaOut => P(8)(524));
U_F9525: entity F port map(lamdaA => P(9)(525),lamdaB => P(9)(527),lamdaOut => P(8)(525));
U_G9526: entity G port map(lamdaA => P(9)(524),lamdaB => P(9)(526),s => s(9)(262),lamdaOut => P(8)(526));
U_G9527: entity G port map(lamdaA => P(9)(525),lamdaB => P(9)(527),s => s(9)(263),lamdaOut => P(8)(527));
U_F9528: entity F port map(lamdaA => P(9)(528),lamdaB => P(9)(530),lamdaOut => P(8)(528));
U_F9529: entity F port map(lamdaA => P(9)(529),lamdaB => P(9)(531),lamdaOut => P(8)(529));
U_G9530: entity G port map(lamdaA => P(9)(528),lamdaB => P(9)(530),s => s(9)(264),lamdaOut => P(8)(530));
U_G9531: entity G port map(lamdaA => P(9)(529),lamdaB => P(9)(531),s => s(9)(265),lamdaOut => P(8)(531));
U_F9532: entity F port map(lamdaA => P(9)(532),lamdaB => P(9)(534),lamdaOut => P(8)(532));
U_F9533: entity F port map(lamdaA => P(9)(533),lamdaB => P(9)(535),lamdaOut => P(8)(533));
U_G9534: entity G port map(lamdaA => P(9)(532),lamdaB => P(9)(534),s => s(9)(266),lamdaOut => P(8)(534));
U_G9535: entity G port map(lamdaA => P(9)(533),lamdaB => P(9)(535),s => s(9)(267),lamdaOut => P(8)(535));
U_F9536: entity F port map(lamdaA => P(9)(536),lamdaB => P(9)(538),lamdaOut => P(8)(536));
U_F9537: entity F port map(lamdaA => P(9)(537),lamdaB => P(9)(539),lamdaOut => P(8)(537));
U_G9538: entity G port map(lamdaA => P(9)(536),lamdaB => P(9)(538),s => s(9)(268),lamdaOut => P(8)(538));
U_G9539: entity G port map(lamdaA => P(9)(537),lamdaB => P(9)(539),s => s(9)(269),lamdaOut => P(8)(539));
U_F9540: entity F port map(lamdaA => P(9)(540),lamdaB => P(9)(542),lamdaOut => P(8)(540));
U_F9541: entity F port map(lamdaA => P(9)(541),lamdaB => P(9)(543),lamdaOut => P(8)(541));
U_G9542: entity G port map(lamdaA => P(9)(540),lamdaB => P(9)(542),s => s(9)(270),lamdaOut => P(8)(542));
U_G9543: entity G port map(lamdaA => P(9)(541),lamdaB => P(9)(543),s => s(9)(271),lamdaOut => P(8)(543));
U_F9544: entity F port map(lamdaA => P(9)(544),lamdaB => P(9)(546),lamdaOut => P(8)(544));
U_F9545: entity F port map(lamdaA => P(9)(545),lamdaB => P(9)(547),lamdaOut => P(8)(545));
U_G9546: entity G port map(lamdaA => P(9)(544),lamdaB => P(9)(546),s => s(9)(272),lamdaOut => P(8)(546));
U_G9547: entity G port map(lamdaA => P(9)(545),lamdaB => P(9)(547),s => s(9)(273),lamdaOut => P(8)(547));
U_F9548: entity F port map(lamdaA => P(9)(548),lamdaB => P(9)(550),lamdaOut => P(8)(548));
U_F9549: entity F port map(lamdaA => P(9)(549),lamdaB => P(9)(551),lamdaOut => P(8)(549));
U_G9550: entity G port map(lamdaA => P(9)(548),lamdaB => P(9)(550),s => s(9)(274),lamdaOut => P(8)(550));
U_G9551: entity G port map(lamdaA => P(9)(549),lamdaB => P(9)(551),s => s(9)(275),lamdaOut => P(8)(551));
U_F9552: entity F port map(lamdaA => P(9)(552),lamdaB => P(9)(554),lamdaOut => P(8)(552));
U_F9553: entity F port map(lamdaA => P(9)(553),lamdaB => P(9)(555),lamdaOut => P(8)(553));
U_G9554: entity G port map(lamdaA => P(9)(552),lamdaB => P(9)(554),s => s(9)(276),lamdaOut => P(8)(554));
U_G9555: entity G port map(lamdaA => P(9)(553),lamdaB => P(9)(555),s => s(9)(277),lamdaOut => P(8)(555));
U_F9556: entity F port map(lamdaA => P(9)(556),lamdaB => P(9)(558),lamdaOut => P(8)(556));
U_F9557: entity F port map(lamdaA => P(9)(557),lamdaB => P(9)(559),lamdaOut => P(8)(557));
U_G9558: entity G port map(lamdaA => P(9)(556),lamdaB => P(9)(558),s => s(9)(278),lamdaOut => P(8)(558));
U_G9559: entity G port map(lamdaA => P(9)(557),lamdaB => P(9)(559),s => s(9)(279),lamdaOut => P(8)(559));
U_F9560: entity F port map(lamdaA => P(9)(560),lamdaB => P(9)(562),lamdaOut => P(8)(560));
U_F9561: entity F port map(lamdaA => P(9)(561),lamdaB => P(9)(563),lamdaOut => P(8)(561));
U_G9562: entity G port map(lamdaA => P(9)(560),lamdaB => P(9)(562),s => s(9)(280),lamdaOut => P(8)(562));
U_G9563: entity G port map(lamdaA => P(9)(561),lamdaB => P(9)(563),s => s(9)(281),lamdaOut => P(8)(563));
U_F9564: entity F port map(lamdaA => P(9)(564),lamdaB => P(9)(566),lamdaOut => P(8)(564));
U_F9565: entity F port map(lamdaA => P(9)(565),lamdaB => P(9)(567),lamdaOut => P(8)(565));
U_G9566: entity G port map(lamdaA => P(9)(564),lamdaB => P(9)(566),s => s(9)(282),lamdaOut => P(8)(566));
U_G9567: entity G port map(lamdaA => P(9)(565),lamdaB => P(9)(567),s => s(9)(283),lamdaOut => P(8)(567));
U_F9568: entity F port map(lamdaA => P(9)(568),lamdaB => P(9)(570),lamdaOut => P(8)(568));
U_F9569: entity F port map(lamdaA => P(9)(569),lamdaB => P(9)(571),lamdaOut => P(8)(569));
U_G9570: entity G port map(lamdaA => P(9)(568),lamdaB => P(9)(570),s => s(9)(284),lamdaOut => P(8)(570));
U_G9571: entity G port map(lamdaA => P(9)(569),lamdaB => P(9)(571),s => s(9)(285),lamdaOut => P(8)(571));
U_F9572: entity F port map(lamdaA => P(9)(572),lamdaB => P(9)(574),lamdaOut => P(8)(572));
U_F9573: entity F port map(lamdaA => P(9)(573),lamdaB => P(9)(575),lamdaOut => P(8)(573));
U_G9574: entity G port map(lamdaA => P(9)(572),lamdaB => P(9)(574),s => s(9)(286),lamdaOut => P(8)(574));
U_G9575: entity G port map(lamdaA => P(9)(573),lamdaB => P(9)(575),s => s(9)(287),lamdaOut => P(8)(575));
U_F9576: entity F port map(lamdaA => P(9)(576),lamdaB => P(9)(578),lamdaOut => P(8)(576));
U_F9577: entity F port map(lamdaA => P(9)(577),lamdaB => P(9)(579),lamdaOut => P(8)(577));
U_G9578: entity G port map(lamdaA => P(9)(576),lamdaB => P(9)(578),s => s(9)(288),lamdaOut => P(8)(578));
U_G9579: entity G port map(lamdaA => P(9)(577),lamdaB => P(9)(579),s => s(9)(289),lamdaOut => P(8)(579));
U_F9580: entity F port map(lamdaA => P(9)(580),lamdaB => P(9)(582),lamdaOut => P(8)(580));
U_F9581: entity F port map(lamdaA => P(9)(581),lamdaB => P(9)(583),lamdaOut => P(8)(581));
U_G9582: entity G port map(lamdaA => P(9)(580),lamdaB => P(9)(582),s => s(9)(290),lamdaOut => P(8)(582));
U_G9583: entity G port map(lamdaA => P(9)(581),lamdaB => P(9)(583),s => s(9)(291),lamdaOut => P(8)(583));
U_F9584: entity F port map(lamdaA => P(9)(584),lamdaB => P(9)(586),lamdaOut => P(8)(584));
U_F9585: entity F port map(lamdaA => P(9)(585),lamdaB => P(9)(587),lamdaOut => P(8)(585));
U_G9586: entity G port map(lamdaA => P(9)(584),lamdaB => P(9)(586),s => s(9)(292),lamdaOut => P(8)(586));
U_G9587: entity G port map(lamdaA => P(9)(585),lamdaB => P(9)(587),s => s(9)(293),lamdaOut => P(8)(587));
U_F9588: entity F port map(lamdaA => P(9)(588),lamdaB => P(9)(590),lamdaOut => P(8)(588));
U_F9589: entity F port map(lamdaA => P(9)(589),lamdaB => P(9)(591),lamdaOut => P(8)(589));
U_G9590: entity G port map(lamdaA => P(9)(588),lamdaB => P(9)(590),s => s(9)(294),lamdaOut => P(8)(590));
U_G9591: entity G port map(lamdaA => P(9)(589),lamdaB => P(9)(591),s => s(9)(295),lamdaOut => P(8)(591));
U_F9592: entity F port map(lamdaA => P(9)(592),lamdaB => P(9)(594),lamdaOut => P(8)(592));
U_F9593: entity F port map(lamdaA => P(9)(593),lamdaB => P(9)(595),lamdaOut => P(8)(593));
U_G9594: entity G port map(lamdaA => P(9)(592),lamdaB => P(9)(594),s => s(9)(296),lamdaOut => P(8)(594));
U_G9595: entity G port map(lamdaA => P(9)(593),lamdaB => P(9)(595),s => s(9)(297),lamdaOut => P(8)(595));
U_F9596: entity F port map(lamdaA => P(9)(596),lamdaB => P(9)(598),lamdaOut => P(8)(596));
U_F9597: entity F port map(lamdaA => P(9)(597),lamdaB => P(9)(599),lamdaOut => P(8)(597));
U_G9598: entity G port map(lamdaA => P(9)(596),lamdaB => P(9)(598),s => s(9)(298),lamdaOut => P(8)(598));
U_G9599: entity G port map(lamdaA => P(9)(597),lamdaB => P(9)(599),s => s(9)(299),lamdaOut => P(8)(599));
U_F9600: entity F port map(lamdaA => P(9)(600),lamdaB => P(9)(602),lamdaOut => P(8)(600));
U_F9601: entity F port map(lamdaA => P(9)(601),lamdaB => P(9)(603),lamdaOut => P(8)(601));
U_G9602: entity G port map(lamdaA => P(9)(600),lamdaB => P(9)(602),s => s(9)(300),lamdaOut => P(8)(602));
U_G9603: entity G port map(lamdaA => P(9)(601),lamdaB => P(9)(603),s => s(9)(301),lamdaOut => P(8)(603));
U_F9604: entity F port map(lamdaA => P(9)(604),lamdaB => P(9)(606),lamdaOut => P(8)(604));
U_F9605: entity F port map(lamdaA => P(9)(605),lamdaB => P(9)(607),lamdaOut => P(8)(605));
U_G9606: entity G port map(lamdaA => P(9)(604),lamdaB => P(9)(606),s => s(9)(302),lamdaOut => P(8)(606));
U_G9607: entity G port map(lamdaA => P(9)(605),lamdaB => P(9)(607),s => s(9)(303),lamdaOut => P(8)(607));
U_F9608: entity F port map(lamdaA => P(9)(608),lamdaB => P(9)(610),lamdaOut => P(8)(608));
U_F9609: entity F port map(lamdaA => P(9)(609),lamdaB => P(9)(611),lamdaOut => P(8)(609));
U_G9610: entity G port map(lamdaA => P(9)(608),lamdaB => P(9)(610),s => s(9)(304),lamdaOut => P(8)(610));
U_G9611: entity G port map(lamdaA => P(9)(609),lamdaB => P(9)(611),s => s(9)(305),lamdaOut => P(8)(611));
U_F9612: entity F port map(lamdaA => P(9)(612),lamdaB => P(9)(614),lamdaOut => P(8)(612));
U_F9613: entity F port map(lamdaA => P(9)(613),lamdaB => P(9)(615),lamdaOut => P(8)(613));
U_G9614: entity G port map(lamdaA => P(9)(612),lamdaB => P(9)(614),s => s(9)(306),lamdaOut => P(8)(614));
U_G9615: entity G port map(lamdaA => P(9)(613),lamdaB => P(9)(615),s => s(9)(307),lamdaOut => P(8)(615));
U_F9616: entity F port map(lamdaA => P(9)(616),lamdaB => P(9)(618),lamdaOut => P(8)(616));
U_F9617: entity F port map(lamdaA => P(9)(617),lamdaB => P(9)(619),lamdaOut => P(8)(617));
U_G9618: entity G port map(lamdaA => P(9)(616),lamdaB => P(9)(618),s => s(9)(308),lamdaOut => P(8)(618));
U_G9619: entity G port map(lamdaA => P(9)(617),lamdaB => P(9)(619),s => s(9)(309),lamdaOut => P(8)(619));
U_F9620: entity F port map(lamdaA => P(9)(620),lamdaB => P(9)(622),lamdaOut => P(8)(620));
U_F9621: entity F port map(lamdaA => P(9)(621),lamdaB => P(9)(623),lamdaOut => P(8)(621));
U_G9622: entity G port map(lamdaA => P(9)(620),lamdaB => P(9)(622),s => s(9)(310),lamdaOut => P(8)(622));
U_G9623: entity G port map(lamdaA => P(9)(621),lamdaB => P(9)(623),s => s(9)(311),lamdaOut => P(8)(623));
U_F9624: entity F port map(lamdaA => P(9)(624),lamdaB => P(9)(626),lamdaOut => P(8)(624));
U_F9625: entity F port map(lamdaA => P(9)(625),lamdaB => P(9)(627),lamdaOut => P(8)(625));
U_G9626: entity G port map(lamdaA => P(9)(624),lamdaB => P(9)(626),s => s(9)(312),lamdaOut => P(8)(626));
U_G9627: entity G port map(lamdaA => P(9)(625),lamdaB => P(9)(627),s => s(9)(313),lamdaOut => P(8)(627));
U_F9628: entity F port map(lamdaA => P(9)(628),lamdaB => P(9)(630),lamdaOut => P(8)(628));
U_F9629: entity F port map(lamdaA => P(9)(629),lamdaB => P(9)(631),lamdaOut => P(8)(629));
U_G9630: entity G port map(lamdaA => P(9)(628),lamdaB => P(9)(630),s => s(9)(314),lamdaOut => P(8)(630));
U_G9631: entity G port map(lamdaA => P(9)(629),lamdaB => P(9)(631),s => s(9)(315),lamdaOut => P(8)(631));
U_F9632: entity F port map(lamdaA => P(9)(632),lamdaB => P(9)(634),lamdaOut => P(8)(632));
U_F9633: entity F port map(lamdaA => P(9)(633),lamdaB => P(9)(635),lamdaOut => P(8)(633));
U_G9634: entity G port map(lamdaA => P(9)(632),lamdaB => P(9)(634),s => s(9)(316),lamdaOut => P(8)(634));
U_G9635: entity G port map(lamdaA => P(9)(633),lamdaB => P(9)(635),s => s(9)(317),lamdaOut => P(8)(635));
U_F9636: entity F port map(lamdaA => P(9)(636),lamdaB => P(9)(638),lamdaOut => P(8)(636));
U_F9637: entity F port map(lamdaA => P(9)(637),lamdaB => P(9)(639),lamdaOut => P(8)(637));
U_G9638: entity G port map(lamdaA => P(9)(636),lamdaB => P(9)(638),s => s(9)(318),lamdaOut => P(8)(638));
U_G9639: entity G port map(lamdaA => P(9)(637),lamdaB => P(9)(639),s => s(9)(319),lamdaOut => P(8)(639));
U_F9640: entity F port map(lamdaA => P(9)(640),lamdaB => P(9)(642),lamdaOut => P(8)(640));
U_F9641: entity F port map(lamdaA => P(9)(641),lamdaB => P(9)(643),lamdaOut => P(8)(641));
U_G9642: entity G port map(lamdaA => P(9)(640),lamdaB => P(9)(642),s => s(9)(320),lamdaOut => P(8)(642));
U_G9643: entity G port map(lamdaA => P(9)(641),lamdaB => P(9)(643),s => s(9)(321),lamdaOut => P(8)(643));
U_F9644: entity F port map(lamdaA => P(9)(644),lamdaB => P(9)(646),lamdaOut => P(8)(644));
U_F9645: entity F port map(lamdaA => P(9)(645),lamdaB => P(9)(647),lamdaOut => P(8)(645));
U_G9646: entity G port map(lamdaA => P(9)(644),lamdaB => P(9)(646),s => s(9)(322),lamdaOut => P(8)(646));
U_G9647: entity G port map(lamdaA => P(9)(645),lamdaB => P(9)(647),s => s(9)(323),lamdaOut => P(8)(647));
U_F9648: entity F port map(lamdaA => P(9)(648),lamdaB => P(9)(650),lamdaOut => P(8)(648));
U_F9649: entity F port map(lamdaA => P(9)(649),lamdaB => P(9)(651),lamdaOut => P(8)(649));
U_G9650: entity G port map(lamdaA => P(9)(648),lamdaB => P(9)(650),s => s(9)(324),lamdaOut => P(8)(650));
U_G9651: entity G port map(lamdaA => P(9)(649),lamdaB => P(9)(651),s => s(9)(325),lamdaOut => P(8)(651));
U_F9652: entity F port map(lamdaA => P(9)(652),lamdaB => P(9)(654),lamdaOut => P(8)(652));
U_F9653: entity F port map(lamdaA => P(9)(653),lamdaB => P(9)(655),lamdaOut => P(8)(653));
U_G9654: entity G port map(lamdaA => P(9)(652),lamdaB => P(9)(654),s => s(9)(326),lamdaOut => P(8)(654));
U_G9655: entity G port map(lamdaA => P(9)(653),lamdaB => P(9)(655),s => s(9)(327),lamdaOut => P(8)(655));
U_F9656: entity F port map(lamdaA => P(9)(656),lamdaB => P(9)(658),lamdaOut => P(8)(656));
U_F9657: entity F port map(lamdaA => P(9)(657),lamdaB => P(9)(659),lamdaOut => P(8)(657));
U_G9658: entity G port map(lamdaA => P(9)(656),lamdaB => P(9)(658),s => s(9)(328),lamdaOut => P(8)(658));
U_G9659: entity G port map(lamdaA => P(9)(657),lamdaB => P(9)(659),s => s(9)(329),lamdaOut => P(8)(659));
U_F9660: entity F port map(lamdaA => P(9)(660),lamdaB => P(9)(662),lamdaOut => P(8)(660));
U_F9661: entity F port map(lamdaA => P(9)(661),lamdaB => P(9)(663),lamdaOut => P(8)(661));
U_G9662: entity G port map(lamdaA => P(9)(660),lamdaB => P(9)(662),s => s(9)(330),lamdaOut => P(8)(662));
U_G9663: entity G port map(lamdaA => P(9)(661),lamdaB => P(9)(663),s => s(9)(331),lamdaOut => P(8)(663));
U_F9664: entity F port map(lamdaA => P(9)(664),lamdaB => P(9)(666),lamdaOut => P(8)(664));
U_F9665: entity F port map(lamdaA => P(9)(665),lamdaB => P(9)(667),lamdaOut => P(8)(665));
U_G9666: entity G port map(lamdaA => P(9)(664),lamdaB => P(9)(666),s => s(9)(332),lamdaOut => P(8)(666));
U_G9667: entity G port map(lamdaA => P(9)(665),lamdaB => P(9)(667),s => s(9)(333),lamdaOut => P(8)(667));
U_F9668: entity F port map(lamdaA => P(9)(668),lamdaB => P(9)(670),lamdaOut => P(8)(668));
U_F9669: entity F port map(lamdaA => P(9)(669),lamdaB => P(9)(671),lamdaOut => P(8)(669));
U_G9670: entity G port map(lamdaA => P(9)(668),lamdaB => P(9)(670),s => s(9)(334),lamdaOut => P(8)(670));
U_G9671: entity G port map(lamdaA => P(9)(669),lamdaB => P(9)(671),s => s(9)(335),lamdaOut => P(8)(671));
U_F9672: entity F port map(lamdaA => P(9)(672),lamdaB => P(9)(674),lamdaOut => P(8)(672));
U_F9673: entity F port map(lamdaA => P(9)(673),lamdaB => P(9)(675),lamdaOut => P(8)(673));
U_G9674: entity G port map(lamdaA => P(9)(672),lamdaB => P(9)(674),s => s(9)(336),lamdaOut => P(8)(674));
U_G9675: entity G port map(lamdaA => P(9)(673),lamdaB => P(9)(675),s => s(9)(337),lamdaOut => P(8)(675));
U_F9676: entity F port map(lamdaA => P(9)(676),lamdaB => P(9)(678),lamdaOut => P(8)(676));
U_F9677: entity F port map(lamdaA => P(9)(677),lamdaB => P(9)(679),lamdaOut => P(8)(677));
U_G9678: entity G port map(lamdaA => P(9)(676),lamdaB => P(9)(678),s => s(9)(338),lamdaOut => P(8)(678));
U_G9679: entity G port map(lamdaA => P(9)(677),lamdaB => P(9)(679),s => s(9)(339),lamdaOut => P(8)(679));
U_F9680: entity F port map(lamdaA => P(9)(680),lamdaB => P(9)(682),lamdaOut => P(8)(680));
U_F9681: entity F port map(lamdaA => P(9)(681),lamdaB => P(9)(683),lamdaOut => P(8)(681));
U_G9682: entity G port map(lamdaA => P(9)(680),lamdaB => P(9)(682),s => s(9)(340),lamdaOut => P(8)(682));
U_G9683: entity G port map(lamdaA => P(9)(681),lamdaB => P(9)(683),s => s(9)(341),lamdaOut => P(8)(683));
U_F9684: entity F port map(lamdaA => P(9)(684),lamdaB => P(9)(686),lamdaOut => P(8)(684));
U_F9685: entity F port map(lamdaA => P(9)(685),lamdaB => P(9)(687),lamdaOut => P(8)(685));
U_G9686: entity G port map(lamdaA => P(9)(684),lamdaB => P(9)(686),s => s(9)(342),lamdaOut => P(8)(686));
U_G9687: entity G port map(lamdaA => P(9)(685),lamdaB => P(9)(687),s => s(9)(343),lamdaOut => P(8)(687));
U_F9688: entity F port map(lamdaA => P(9)(688),lamdaB => P(9)(690),lamdaOut => P(8)(688));
U_F9689: entity F port map(lamdaA => P(9)(689),lamdaB => P(9)(691),lamdaOut => P(8)(689));
U_G9690: entity G port map(lamdaA => P(9)(688),lamdaB => P(9)(690),s => s(9)(344),lamdaOut => P(8)(690));
U_G9691: entity G port map(lamdaA => P(9)(689),lamdaB => P(9)(691),s => s(9)(345),lamdaOut => P(8)(691));
U_F9692: entity F port map(lamdaA => P(9)(692),lamdaB => P(9)(694),lamdaOut => P(8)(692));
U_F9693: entity F port map(lamdaA => P(9)(693),lamdaB => P(9)(695),lamdaOut => P(8)(693));
U_G9694: entity G port map(lamdaA => P(9)(692),lamdaB => P(9)(694),s => s(9)(346),lamdaOut => P(8)(694));
U_G9695: entity G port map(lamdaA => P(9)(693),lamdaB => P(9)(695),s => s(9)(347),lamdaOut => P(8)(695));
U_F9696: entity F port map(lamdaA => P(9)(696),lamdaB => P(9)(698),lamdaOut => P(8)(696));
U_F9697: entity F port map(lamdaA => P(9)(697),lamdaB => P(9)(699),lamdaOut => P(8)(697));
U_G9698: entity G port map(lamdaA => P(9)(696),lamdaB => P(9)(698),s => s(9)(348),lamdaOut => P(8)(698));
U_G9699: entity G port map(lamdaA => P(9)(697),lamdaB => P(9)(699),s => s(9)(349),lamdaOut => P(8)(699));
U_F9700: entity F port map(lamdaA => P(9)(700),lamdaB => P(9)(702),lamdaOut => P(8)(700));
U_F9701: entity F port map(lamdaA => P(9)(701),lamdaB => P(9)(703),lamdaOut => P(8)(701));
U_G9702: entity G port map(lamdaA => P(9)(700),lamdaB => P(9)(702),s => s(9)(350),lamdaOut => P(8)(702));
U_G9703: entity G port map(lamdaA => P(9)(701),lamdaB => P(9)(703),s => s(9)(351),lamdaOut => P(8)(703));
U_F9704: entity F port map(lamdaA => P(9)(704),lamdaB => P(9)(706),lamdaOut => P(8)(704));
U_F9705: entity F port map(lamdaA => P(9)(705),lamdaB => P(9)(707),lamdaOut => P(8)(705));
U_G9706: entity G port map(lamdaA => P(9)(704),lamdaB => P(9)(706),s => s(9)(352),lamdaOut => P(8)(706));
U_G9707: entity G port map(lamdaA => P(9)(705),lamdaB => P(9)(707),s => s(9)(353),lamdaOut => P(8)(707));
U_F9708: entity F port map(lamdaA => P(9)(708),lamdaB => P(9)(710),lamdaOut => P(8)(708));
U_F9709: entity F port map(lamdaA => P(9)(709),lamdaB => P(9)(711),lamdaOut => P(8)(709));
U_G9710: entity G port map(lamdaA => P(9)(708),lamdaB => P(9)(710),s => s(9)(354),lamdaOut => P(8)(710));
U_G9711: entity G port map(lamdaA => P(9)(709),lamdaB => P(9)(711),s => s(9)(355),lamdaOut => P(8)(711));
U_F9712: entity F port map(lamdaA => P(9)(712),lamdaB => P(9)(714),lamdaOut => P(8)(712));
U_F9713: entity F port map(lamdaA => P(9)(713),lamdaB => P(9)(715),lamdaOut => P(8)(713));
U_G9714: entity G port map(lamdaA => P(9)(712),lamdaB => P(9)(714),s => s(9)(356),lamdaOut => P(8)(714));
U_G9715: entity G port map(lamdaA => P(9)(713),lamdaB => P(9)(715),s => s(9)(357),lamdaOut => P(8)(715));
U_F9716: entity F port map(lamdaA => P(9)(716),lamdaB => P(9)(718),lamdaOut => P(8)(716));
U_F9717: entity F port map(lamdaA => P(9)(717),lamdaB => P(9)(719),lamdaOut => P(8)(717));
U_G9718: entity G port map(lamdaA => P(9)(716),lamdaB => P(9)(718),s => s(9)(358),lamdaOut => P(8)(718));
U_G9719: entity G port map(lamdaA => P(9)(717),lamdaB => P(9)(719),s => s(9)(359),lamdaOut => P(8)(719));
U_F9720: entity F port map(lamdaA => P(9)(720),lamdaB => P(9)(722),lamdaOut => P(8)(720));
U_F9721: entity F port map(lamdaA => P(9)(721),lamdaB => P(9)(723),lamdaOut => P(8)(721));
U_G9722: entity G port map(lamdaA => P(9)(720),lamdaB => P(9)(722),s => s(9)(360),lamdaOut => P(8)(722));
U_G9723: entity G port map(lamdaA => P(9)(721),lamdaB => P(9)(723),s => s(9)(361),lamdaOut => P(8)(723));
U_F9724: entity F port map(lamdaA => P(9)(724),lamdaB => P(9)(726),lamdaOut => P(8)(724));
U_F9725: entity F port map(lamdaA => P(9)(725),lamdaB => P(9)(727),lamdaOut => P(8)(725));
U_G9726: entity G port map(lamdaA => P(9)(724),lamdaB => P(9)(726),s => s(9)(362),lamdaOut => P(8)(726));
U_G9727: entity G port map(lamdaA => P(9)(725),lamdaB => P(9)(727),s => s(9)(363),lamdaOut => P(8)(727));
U_F9728: entity F port map(lamdaA => P(9)(728),lamdaB => P(9)(730),lamdaOut => P(8)(728));
U_F9729: entity F port map(lamdaA => P(9)(729),lamdaB => P(9)(731),lamdaOut => P(8)(729));
U_G9730: entity G port map(lamdaA => P(9)(728),lamdaB => P(9)(730),s => s(9)(364),lamdaOut => P(8)(730));
U_G9731: entity G port map(lamdaA => P(9)(729),lamdaB => P(9)(731),s => s(9)(365),lamdaOut => P(8)(731));
U_F9732: entity F port map(lamdaA => P(9)(732),lamdaB => P(9)(734),lamdaOut => P(8)(732));
U_F9733: entity F port map(lamdaA => P(9)(733),lamdaB => P(9)(735),lamdaOut => P(8)(733));
U_G9734: entity G port map(lamdaA => P(9)(732),lamdaB => P(9)(734),s => s(9)(366),lamdaOut => P(8)(734));
U_G9735: entity G port map(lamdaA => P(9)(733),lamdaB => P(9)(735),s => s(9)(367),lamdaOut => P(8)(735));
U_F9736: entity F port map(lamdaA => P(9)(736),lamdaB => P(9)(738),lamdaOut => P(8)(736));
U_F9737: entity F port map(lamdaA => P(9)(737),lamdaB => P(9)(739),lamdaOut => P(8)(737));
U_G9738: entity G port map(lamdaA => P(9)(736),lamdaB => P(9)(738),s => s(9)(368),lamdaOut => P(8)(738));
U_G9739: entity G port map(lamdaA => P(9)(737),lamdaB => P(9)(739),s => s(9)(369),lamdaOut => P(8)(739));
U_F9740: entity F port map(lamdaA => P(9)(740),lamdaB => P(9)(742),lamdaOut => P(8)(740));
U_F9741: entity F port map(lamdaA => P(9)(741),lamdaB => P(9)(743),lamdaOut => P(8)(741));
U_G9742: entity G port map(lamdaA => P(9)(740),lamdaB => P(9)(742),s => s(9)(370),lamdaOut => P(8)(742));
U_G9743: entity G port map(lamdaA => P(9)(741),lamdaB => P(9)(743),s => s(9)(371),lamdaOut => P(8)(743));
U_F9744: entity F port map(lamdaA => P(9)(744),lamdaB => P(9)(746),lamdaOut => P(8)(744));
U_F9745: entity F port map(lamdaA => P(9)(745),lamdaB => P(9)(747),lamdaOut => P(8)(745));
U_G9746: entity G port map(lamdaA => P(9)(744),lamdaB => P(9)(746),s => s(9)(372),lamdaOut => P(8)(746));
U_G9747: entity G port map(lamdaA => P(9)(745),lamdaB => P(9)(747),s => s(9)(373),lamdaOut => P(8)(747));
U_F9748: entity F port map(lamdaA => P(9)(748),lamdaB => P(9)(750),lamdaOut => P(8)(748));
U_F9749: entity F port map(lamdaA => P(9)(749),lamdaB => P(9)(751),lamdaOut => P(8)(749));
U_G9750: entity G port map(lamdaA => P(9)(748),lamdaB => P(9)(750),s => s(9)(374),lamdaOut => P(8)(750));
U_G9751: entity G port map(lamdaA => P(9)(749),lamdaB => P(9)(751),s => s(9)(375),lamdaOut => P(8)(751));
U_F9752: entity F port map(lamdaA => P(9)(752),lamdaB => P(9)(754),lamdaOut => P(8)(752));
U_F9753: entity F port map(lamdaA => P(9)(753),lamdaB => P(9)(755),lamdaOut => P(8)(753));
U_G9754: entity G port map(lamdaA => P(9)(752),lamdaB => P(9)(754),s => s(9)(376),lamdaOut => P(8)(754));
U_G9755: entity G port map(lamdaA => P(9)(753),lamdaB => P(9)(755),s => s(9)(377),lamdaOut => P(8)(755));
U_F9756: entity F port map(lamdaA => P(9)(756),lamdaB => P(9)(758),lamdaOut => P(8)(756));
U_F9757: entity F port map(lamdaA => P(9)(757),lamdaB => P(9)(759),lamdaOut => P(8)(757));
U_G9758: entity G port map(lamdaA => P(9)(756),lamdaB => P(9)(758),s => s(9)(378),lamdaOut => P(8)(758));
U_G9759: entity G port map(lamdaA => P(9)(757),lamdaB => P(9)(759),s => s(9)(379),lamdaOut => P(8)(759));
U_F9760: entity F port map(lamdaA => P(9)(760),lamdaB => P(9)(762),lamdaOut => P(8)(760));
U_F9761: entity F port map(lamdaA => P(9)(761),lamdaB => P(9)(763),lamdaOut => P(8)(761));
U_G9762: entity G port map(lamdaA => P(9)(760),lamdaB => P(9)(762),s => s(9)(380),lamdaOut => P(8)(762));
U_G9763: entity G port map(lamdaA => P(9)(761),lamdaB => P(9)(763),s => s(9)(381),lamdaOut => P(8)(763));
U_F9764: entity F port map(lamdaA => P(9)(764),lamdaB => P(9)(766),lamdaOut => P(8)(764));
U_F9765: entity F port map(lamdaA => P(9)(765),lamdaB => P(9)(767),lamdaOut => P(8)(765));
U_G9766: entity G port map(lamdaA => P(9)(764),lamdaB => P(9)(766),s => s(9)(382),lamdaOut => P(8)(766));
U_G9767: entity G port map(lamdaA => P(9)(765),lamdaB => P(9)(767),s => s(9)(383),lamdaOut => P(8)(767));
U_F9768: entity F port map(lamdaA => P(9)(768),lamdaB => P(9)(770),lamdaOut => P(8)(768));
U_F9769: entity F port map(lamdaA => P(9)(769),lamdaB => P(9)(771),lamdaOut => P(8)(769));
U_G9770: entity G port map(lamdaA => P(9)(768),lamdaB => P(9)(770),s => s(9)(384),lamdaOut => P(8)(770));
U_G9771: entity G port map(lamdaA => P(9)(769),lamdaB => P(9)(771),s => s(9)(385),lamdaOut => P(8)(771));
U_F9772: entity F port map(lamdaA => P(9)(772),lamdaB => P(9)(774),lamdaOut => P(8)(772));
U_F9773: entity F port map(lamdaA => P(9)(773),lamdaB => P(9)(775),lamdaOut => P(8)(773));
U_G9774: entity G port map(lamdaA => P(9)(772),lamdaB => P(9)(774),s => s(9)(386),lamdaOut => P(8)(774));
U_G9775: entity G port map(lamdaA => P(9)(773),lamdaB => P(9)(775),s => s(9)(387),lamdaOut => P(8)(775));
U_F9776: entity F port map(lamdaA => P(9)(776),lamdaB => P(9)(778),lamdaOut => P(8)(776));
U_F9777: entity F port map(lamdaA => P(9)(777),lamdaB => P(9)(779),lamdaOut => P(8)(777));
U_G9778: entity G port map(lamdaA => P(9)(776),lamdaB => P(9)(778),s => s(9)(388),lamdaOut => P(8)(778));
U_G9779: entity G port map(lamdaA => P(9)(777),lamdaB => P(9)(779),s => s(9)(389),lamdaOut => P(8)(779));
U_F9780: entity F port map(lamdaA => P(9)(780),lamdaB => P(9)(782),lamdaOut => P(8)(780));
U_F9781: entity F port map(lamdaA => P(9)(781),lamdaB => P(9)(783),lamdaOut => P(8)(781));
U_G9782: entity G port map(lamdaA => P(9)(780),lamdaB => P(9)(782),s => s(9)(390),lamdaOut => P(8)(782));
U_G9783: entity G port map(lamdaA => P(9)(781),lamdaB => P(9)(783),s => s(9)(391),lamdaOut => P(8)(783));
U_F9784: entity F port map(lamdaA => P(9)(784),lamdaB => P(9)(786),lamdaOut => P(8)(784));
U_F9785: entity F port map(lamdaA => P(9)(785),lamdaB => P(9)(787),lamdaOut => P(8)(785));
U_G9786: entity G port map(lamdaA => P(9)(784),lamdaB => P(9)(786),s => s(9)(392),lamdaOut => P(8)(786));
U_G9787: entity G port map(lamdaA => P(9)(785),lamdaB => P(9)(787),s => s(9)(393),lamdaOut => P(8)(787));
U_F9788: entity F port map(lamdaA => P(9)(788),lamdaB => P(9)(790),lamdaOut => P(8)(788));
U_F9789: entity F port map(lamdaA => P(9)(789),lamdaB => P(9)(791),lamdaOut => P(8)(789));
U_G9790: entity G port map(lamdaA => P(9)(788),lamdaB => P(9)(790),s => s(9)(394),lamdaOut => P(8)(790));
U_G9791: entity G port map(lamdaA => P(9)(789),lamdaB => P(9)(791),s => s(9)(395),lamdaOut => P(8)(791));
U_F9792: entity F port map(lamdaA => P(9)(792),lamdaB => P(9)(794),lamdaOut => P(8)(792));
U_F9793: entity F port map(lamdaA => P(9)(793),lamdaB => P(9)(795),lamdaOut => P(8)(793));
U_G9794: entity G port map(lamdaA => P(9)(792),lamdaB => P(9)(794),s => s(9)(396),lamdaOut => P(8)(794));
U_G9795: entity G port map(lamdaA => P(9)(793),lamdaB => P(9)(795),s => s(9)(397),lamdaOut => P(8)(795));
U_F9796: entity F port map(lamdaA => P(9)(796),lamdaB => P(9)(798),lamdaOut => P(8)(796));
U_F9797: entity F port map(lamdaA => P(9)(797),lamdaB => P(9)(799),lamdaOut => P(8)(797));
U_G9798: entity G port map(lamdaA => P(9)(796),lamdaB => P(9)(798),s => s(9)(398),lamdaOut => P(8)(798));
U_G9799: entity G port map(lamdaA => P(9)(797),lamdaB => P(9)(799),s => s(9)(399),lamdaOut => P(8)(799));
U_F9800: entity F port map(lamdaA => P(9)(800),lamdaB => P(9)(802),lamdaOut => P(8)(800));
U_F9801: entity F port map(lamdaA => P(9)(801),lamdaB => P(9)(803),lamdaOut => P(8)(801));
U_G9802: entity G port map(lamdaA => P(9)(800),lamdaB => P(9)(802),s => s(9)(400),lamdaOut => P(8)(802));
U_G9803: entity G port map(lamdaA => P(9)(801),lamdaB => P(9)(803),s => s(9)(401),lamdaOut => P(8)(803));
U_F9804: entity F port map(lamdaA => P(9)(804),lamdaB => P(9)(806),lamdaOut => P(8)(804));
U_F9805: entity F port map(lamdaA => P(9)(805),lamdaB => P(9)(807),lamdaOut => P(8)(805));
U_G9806: entity G port map(lamdaA => P(9)(804),lamdaB => P(9)(806),s => s(9)(402),lamdaOut => P(8)(806));
U_G9807: entity G port map(lamdaA => P(9)(805),lamdaB => P(9)(807),s => s(9)(403),lamdaOut => P(8)(807));
U_F9808: entity F port map(lamdaA => P(9)(808),lamdaB => P(9)(810),lamdaOut => P(8)(808));
U_F9809: entity F port map(lamdaA => P(9)(809),lamdaB => P(9)(811),lamdaOut => P(8)(809));
U_G9810: entity G port map(lamdaA => P(9)(808),lamdaB => P(9)(810),s => s(9)(404),lamdaOut => P(8)(810));
U_G9811: entity G port map(lamdaA => P(9)(809),lamdaB => P(9)(811),s => s(9)(405),lamdaOut => P(8)(811));
U_F9812: entity F port map(lamdaA => P(9)(812),lamdaB => P(9)(814),lamdaOut => P(8)(812));
U_F9813: entity F port map(lamdaA => P(9)(813),lamdaB => P(9)(815),lamdaOut => P(8)(813));
U_G9814: entity G port map(lamdaA => P(9)(812),lamdaB => P(9)(814),s => s(9)(406),lamdaOut => P(8)(814));
U_G9815: entity G port map(lamdaA => P(9)(813),lamdaB => P(9)(815),s => s(9)(407),lamdaOut => P(8)(815));
U_F9816: entity F port map(lamdaA => P(9)(816),lamdaB => P(9)(818),lamdaOut => P(8)(816));
U_F9817: entity F port map(lamdaA => P(9)(817),lamdaB => P(9)(819),lamdaOut => P(8)(817));
U_G9818: entity G port map(lamdaA => P(9)(816),lamdaB => P(9)(818),s => s(9)(408),lamdaOut => P(8)(818));
U_G9819: entity G port map(lamdaA => P(9)(817),lamdaB => P(9)(819),s => s(9)(409),lamdaOut => P(8)(819));
U_F9820: entity F port map(lamdaA => P(9)(820),lamdaB => P(9)(822),lamdaOut => P(8)(820));
U_F9821: entity F port map(lamdaA => P(9)(821),lamdaB => P(9)(823),lamdaOut => P(8)(821));
U_G9822: entity G port map(lamdaA => P(9)(820),lamdaB => P(9)(822),s => s(9)(410),lamdaOut => P(8)(822));
U_G9823: entity G port map(lamdaA => P(9)(821),lamdaB => P(9)(823),s => s(9)(411),lamdaOut => P(8)(823));
U_F9824: entity F port map(lamdaA => P(9)(824),lamdaB => P(9)(826),lamdaOut => P(8)(824));
U_F9825: entity F port map(lamdaA => P(9)(825),lamdaB => P(9)(827),lamdaOut => P(8)(825));
U_G9826: entity G port map(lamdaA => P(9)(824),lamdaB => P(9)(826),s => s(9)(412),lamdaOut => P(8)(826));
U_G9827: entity G port map(lamdaA => P(9)(825),lamdaB => P(9)(827),s => s(9)(413),lamdaOut => P(8)(827));
U_F9828: entity F port map(lamdaA => P(9)(828),lamdaB => P(9)(830),lamdaOut => P(8)(828));
U_F9829: entity F port map(lamdaA => P(9)(829),lamdaB => P(9)(831),lamdaOut => P(8)(829));
U_G9830: entity G port map(lamdaA => P(9)(828),lamdaB => P(9)(830),s => s(9)(414),lamdaOut => P(8)(830));
U_G9831: entity G port map(lamdaA => P(9)(829),lamdaB => P(9)(831),s => s(9)(415),lamdaOut => P(8)(831));
U_F9832: entity F port map(lamdaA => P(9)(832),lamdaB => P(9)(834),lamdaOut => P(8)(832));
U_F9833: entity F port map(lamdaA => P(9)(833),lamdaB => P(9)(835),lamdaOut => P(8)(833));
U_G9834: entity G port map(lamdaA => P(9)(832),lamdaB => P(9)(834),s => s(9)(416),lamdaOut => P(8)(834));
U_G9835: entity G port map(lamdaA => P(9)(833),lamdaB => P(9)(835),s => s(9)(417),lamdaOut => P(8)(835));
U_F9836: entity F port map(lamdaA => P(9)(836),lamdaB => P(9)(838),lamdaOut => P(8)(836));
U_F9837: entity F port map(lamdaA => P(9)(837),lamdaB => P(9)(839),lamdaOut => P(8)(837));
U_G9838: entity G port map(lamdaA => P(9)(836),lamdaB => P(9)(838),s => s(9)(418),lamdaOut => P(8)(838));
U_G9839: entity G port map(lamdaA => P(9)(837),lamdaB => P(9)(839),s => s(9)(419),lamdaOut => P(8)(839));
U_F9840: entity F port map(lamdaA => P(9)(840),lamdaB => P(9)(842),lamdaOut => P(8)(840));
U_F9841: entity F port map(lamdaA => P(9)(841),lamdaB => P(9)(843),lamdaOut => P(8)(841));
U_G9842: entity G port map(lamdaA => P(9)(840),lamdaB => P(9)(842),s => s(9)(420),lamdaOut => P(8)(842));
U_G9843: entity G port map(lamdaA => P(9)(841),lamdaB => P(9)(843),s => s(9)(421),lamdaOut => P(8)(843));
U_F9844: entity F port map(lamdaA => P(9)(844),lamdaB => P(9)(846),lamdaOut => P(8)(844));
U_F9845: entity F port map(lamdaA => P(9)(845),lamdaB => P(9)(847),lamdaOut => P(8)(845));
U_G9846: entity G port map(lamdaA => P(9)(844),lamdaB => P(9)(846),s => s(9)(422),lamdaOut => P(8)(846));
U_G9847: entity G port map(lamdaA => P(9)(845),lamdaB => P(9)(847),s => s(9)(423),lamdaOut => P(8)(847));
U_F9848: entity F port map(lamdaA => P(9)(848),lamdaB => P(9)(850),lamdaOut => P(8)(848));
U_F9849: entity F port map(lamdaA => P(9)(849),lamdaB => P(9)(851),lamdaOut => P(8)(849));
U_G9850: entity G port map(lamdaA => P(9)(848),lamdaB => P(9)(850),s => s(9)(424),lamdaOut => P(8)(850));
U_G9851: entity G port map(lamdaA => P(9)(849),lamdaB => P(9)(851),s => s(9)(425),lamdaOut => P(8)(851));
U_F9852: entity F port map(lamdaA => P(9)(852),lamdaB => P(9)(854),lamdaOut => P(8)(852));
U_F9853: entity F port map(lamdaA => P(9)(853),lamdaB => P(9)(855),lamdaOut => P(8)(853));
U_G9854: entity G port map(lamdaA => P(9)(852),lamdaB => P(9)(854),s => s(9)(426),lamdaOut => P(8)(854));
U_G9855: entity G port map(lamdaA => P(9)(853),lamdaB => P(9)(855),s => s(9)(427),lamdaOut => P(8)(855));
U_F9856: entity F port map(lamdaA => P(9)(856),lamdaB => P(9)(858),lamdaOut => P(8)(856));
U_F9857: entity F port map(lamdaA => P(9)(857),lamdaB => P(9)(859),lamdaOut => P(8)(857));
U_G9858: entity G port map(lamdaA => P(9)(856),lamdaB => P(9)(858),s => s(9)(428),lamdaOut => P(8)(858));
U_G9859: entity G port map(lamdaA => P(9)(857),lamdaB => P(9)(859),s => s(9)(429),lamdaOut => P(8)(859));
U_F9860: entity F port map(lamdaA => P(9)(860),lamdaB => P(9)(862),lamdaOut => P(8)(860));
U_F9861: entity F port map(lamdaA => P(9)(861),lamdaB => P(9)(863),lamdaOut => P(8)(861));
U_G9862: entity G port map(lamdaA => P(9)(860),lamdaB => P(9)(862),s => s(9)(430),lamdaOut => P(8)(862));
U_G9863: entity G port map(lamdaA => P(9)(861),lamdaB => P(9)(863),s => s(9)(431),lamdaOut => P(8)(863));
U_F9864: entity F port map(lamdaA => P(9)(864),lamdaB => P(9)(866),lamdaOut => P(8)(864));
U_F9865: entity F port map(lamdaA => P(9)(865),lamdaB => P(9)(867),lamdaOut => P(8)(865));
U_G9866: entity G port map(lamdaA => P(9)(864),lamdaB => P(9)(866),s => s(9)(432),lamdaOut => P(8)(866));
U_G9867: entity G port map(lamdaA => P(9)(865),lamdaB => P(9)(867),s => s(9)(433),lamdaOut => P(8)(867));
U_F9868: entity F port map(lamdaA => P(9)(868),lamdaB => P(9)(870),lamdaOut => P(8)(868));
U_F9869: entity F port map(lamdaA => P(9)(869),lamdaB => P(9)(871),lamdaOut => P(8)(869));
U_G9870: entity G port map(lamdaA => P(9)(868),lamdaB => P(9)(870),s => s(9)(434),lamdaOut => P(8)(870));
U_G9871: entity G port map(lamdaA => P(9)(869),lamdaB => P(9)(871),s => s(9)(435),lamdaOut => P(8)(871));
U_F9872: entity F port map(lamdaA => P(9)(872),lamdaB => P(9)(874),lamdaOut => P(8)(872));
U_F9873: entity F port map(lamdaA => P(9)(873),lamdaB => P(9)(875),lamdaOut => P(8)(873));
U_G9874: entity G port map(lamdaA => P(9)(872),lamdaB => P(9)(874),s => s(9)(436),lamdaOut => P(8)(874));
U_G9875: entity G port map(lamdaA => P(9)(873),lamdaB => P(9)(875),s => s(9)(437),lamdaOut => P(8)(875));
U_F9876: entity F port map(lamdaA => P(9)(876),lamdaB => P(9)(878),lamdaOut => P(8)(876));
U_F9877: entity F port map(lamdaA => P(9)(877),lamdaB => P(9)(879),lamdaOut => P(8)(877));
U_G9878: entity G port map(lamdaA => P(9)(876),lamdaB => P(9)(878),s => s(9)(438),lamdaOut => P(8)(878));
U_G9879: entity G port map(lamdaA => P(9)(877),lamdaB => P(9)(879),s => s(9)(439),lamdaOut => P(8)(879));
U_F9880: entity F port map(lamdaA => P(9)(880),lamdaB => P(9)(882),lamdaOut => P(8)(880));
U_F9881: entity F port map(lamdaA => P(9)(881),lamdaB => P(9)(883),lamdaOut => P(8)(881));
U_G9882: entity G port map(lamdaA => P(9)(880),lamdaB => P(9)(882),s => s(9)(440),lamdaOut => P(8)(882));
U_G9883: entity G port map(lamdaA => P(9)(881),lamdaB => P(9)(883),s => s(9)(441),lamdaOut => P(8)(883));
U_F9884: entity F port map(lamdaA => P(9)(884),lamdaB => P(9)(886),lamdaOut => P(8)(884));
U_F9885: entity F port map(lamdaA => P(9)(885),lamdaB => P(9)(887),lamdaOut => P(8)(885));
U_G9886: entity G port map(lamdaA => P(9)(884),lamdaB => P(9)(886),s => s(9)(442),lamdaOut => P(8)(886));
U_G9887: entity G port map(lamdaA => P(9)(885),lamdaB => P(9)(887),s => s(9)(443),lamdaOut => P(8)(887));
U_F9888: entity F port map(lamdaA => P(9)(888),lamdaB => P(9)(890),lamdaOut => P(8)(888));
U_F9889: entity F port map(lamdaA => P(9)(889),lamdaB => P(9)(891),lamdaOut => P(8)(889));
U_G9890: entity G port map(lamdaA => P(9)(888),lamdaB => P(9)(890),s => s(9)(444),lamdaOut => P(8)(890));
U_G9891: entity G port map(lamdaA => P(9)(889),lamdaB => P(9)(891),s => s(9)(445),lamdaOut => P(8)(891));
U_F9892: entity F port map(lamdaA => P(9)(892),lamdaB => P(9)(894),lamdaOut => P(8)(892));
U_F9893: entity F port map(lamdaA => P(9)(893),lamdaB => P(9)(895),lamdaOut => P(8)(893));
U_G9894: entity G port map(lamdaA => P(9)(892),lamdaB => P(9)(894),s => s(9)(446),lamdaOut => P(8)(894));
U_G9895: entity G port map(lamdaA => P(9)(893),lamdaB => P(9)(895),s => s(9)(447),lamdaOut => P(8)(895));
U_F9896: entity F port map(lamdaA => P(9)(896),lamdaB => P(9)(898),lamdaOut => P(8)(896));
U_F9897: entity F port map(lamdaA => P(9)(897),lamdaB => P(9)(899),lamdaOut => P(8)(897));
U_G9898: entity G port map(lamdaA => P(9)(896),lamdaB => P(9)(898),s => s(9)(448),lamdaOut => P(8)(898));
U_G9899: entity G port map(lamdaA => P(9)(897),lamdaB => P(9)(899),s => s(9)(449),lamdaOut => P(8)(899));
U_F9900: entity F port map(lamdaA => P(9)(900),lamdaB => P(9)(902),lamdaOut => P(8)(900));
U_F9901: entity F port map(lamdaA => P(9)(901),lamdaB => P(9)(903),lamdaOut => P(8)(901));
U_G9902: entity G port map(lamdaA => P(9)(900),lamdaB => P(9)(902),s => s(9)(450),lamdaOut => P(8)(902));
U_G9903: entity G port map(lamdaA => P(9)(901),lamdaB => P(9)(903),s => s(9)(451),lamdaOut => P(8)(903));
U_F9904: entity F port map(lamdaA => P(9)(904),lamdaB => P(9)(906),lamdaOut => P(8)(904));
U_F9905: entity F port map(lamdaA => P(9)(905),lamdaB => P(9)(907),lamdaOut => P(8)(905));
U_G9906: entity G port map(lamdaA => P(9)(904),lamdaB => P(9)(906),s => s(9)(452),lamdaOut => P(8)(906));
U_G9907: entity G port map(lamdaA => P(9)(905),lamdaB => P(9)(907),s => s(9)(453),lamdaOut => P(8)(907));
U_F9908: entity F port map(lamdaA => P(9)(908),lamdaB => P(9)(910),lamdaOut => P(8)(908));
U_F9909: entity F port map(lamdaA => P(9)(909),lamdaB => P(9)(911),lamdaOut => P(8)(909));
U_G9910: entity G port map(lamdaA => P(9)(908),lamdaB => P(9)(910),s => s(9)(454),lamdaOut => P(8)(910));
U_G9911: entity G port map(lamdaA => P(9)(909),lamdaB => P(9)(911),s => s(9)(455),lamdaOut => P(8)(911));
U_F9912: entity F port map(lamdaA => P(9)(912),lamdaB => P(9)(914),lamdaOut => P(8)(912));
U_F9913: entity F port map(lamdaA => P(9)(913),lamdaB => P(9)(915),lamdaOut => P(8)(913));
U_G9914: entity G port map(lamdaA => P(9)(912),lamdaB => P(9)(914),s => s(9)(456),lamdaOut => P(8)(914));
U_G9915: entity G port map(lamdaA => P(9)(913),lamdaB => P(9)(915),s => s(9)(457),lamdaOut => P(8)(915));
U_F9916: entity F port map(lamdaA => P(9)(916),lamdaB => P(9)(918),lamdaOut => P(8)(916));
U_F9917: entity F port map(lamdaA => P(9)(917),lamdaB => P(9)(919),lamdaOut => P(8)(917));
U_G9918: entity G port map(lamdaA => P(9)(916),lamdaB => P(9)(918),s => s(9)(458),lamdaOut => P(8)(918));
U_G9919: entity G port map(lamdaA => P(9)(917),lamdaB => P(9)(919),s => s(9)(459),lamdaOut => P(8)(919));
U_F9920: entity F port map(lamdaA => P(9)(920),lamdaB => P(9)(922),lamdaOut => P(8)(920));
U_F9921: entity F port map(lamdaA => P(9)(921),lamdaB => P(9)(923),lamdaOut => P(8)(921));
U_G9922: entity G port map(lamdaA => P(9)(920),lamdaB => P(9)(922),s => s(9)(460),lamdaOut => P(8)(922));
U_G9923: entity G port map(lamdaA => P(9)(921),lamdaB => P(9)(923),s => s(9)(461),lamdaOut => P(8)(923));
U_F9924: entity F port map(lamdaA => P(9)(924),lamdaB => P(9)(926),lamdaOut => P(8)(924));
U_F9925: entity F port map(lamdaA => P(9)(925),lamdaB => P(9)(927),lamdaOut => P(8)(925));
U_G9926: entity G port map(lamdaA => P(9)(924),lamdaB => P(9)(926),s => s(9)(462),lamdaOut => P(8)(926));
U_G9927: entity G port map(lamdaA => P(9)(925),lamdaB => P(9)(927),s => s(9)(463),lamdaOut => P(8)(927));
U_F9928: entity F port map(lamdaA => P(9)(928),lamdaB => P(9)(930),lamdaOut => P(8)(928));
U_F9929: entity F port map(lamdaA => P(9)(929),lamdaB => P(9)(931),lamdaOut => P(8)(929));
U_G9930: entity G port map(lamdaA => P(9)(928),lamdaB => P(9)(930),s => s(9)(464),lamdaOut => P(8)(930));
U_G9931: entity G port map(lamdaA => P(9)(929),lamdaB => P(9)(931),s => s(9)(465),lamdaOut => P(8)(931));
U_F9932: entity F port map(lamdaA => P(9)(932),lamdaB => P(9)(934),lamdaOut => P(8)(932));
U_F9933: entity F port map(lamdaA => P(9)(933),lamdaB => P(9)(935),lamdaOut => P(8)(933));
U_G9934: entity G port map(lamdaA => P(9)(932),lamdaB => P(9)(934),s => s(9)(466),lamdaOut => P(8)(934));
U_G9935: entity G port map(lamdaA => P(9)(933),lamdaB => P(9)(935),s => s(9)(467),lamdaOut => P(8)(935));
U_F9936: entity F port map(lamdaA => P(9)(936),lamdaB => P(9)(938),lamdaOut => P(8)(936));
U_F9937: entity F port map(lamdaA => P(9)(937),lamdaB => P(9)(939),lamdaOut => P(8)(937));
U_G9938: entity G port map(lamdaA => P(9)(936),lamdaB => P(9)(938),s => s(9)(468),lamdaOut => P(8)(938));
U_G9939: entity G port map(lamdaA => P(9)(937),lamdaB => P(9)(939),s => s(9)(469),lamdaOut => P(8)(939));
U_F9940: entity F port map(lamdaA => P(9)(940),lamdaB => P(9)(942),lamdaOut => P(8)(940));
U_F9941: entity F port map(lamdaA => P(9)(941),lamdaB => P(9)(943),lamdaOut => P(8)(941));
U_G9942: entity G port map(lamdaA => P(9)(940),lamdaB => P(9)(942),s => s(9)(470),lamdaOut => P(8)(942));
U_G9943: entity G port map(lamdaA => P(9)(941),lamdaB => P(9)(943),s => s(9)(471),lamdaOut => P(8)(943));
U_F9944: entity F port map(lamdaA => P(9)(944),lamdaB => P(9)(946),lamdaOut => P(8)(944));
U_F9945: entity F port map(lamdaA => P(9)(945),lamdaB => P(9)(947),lamdaOut => P(8)(945));
U_G9946: entity G port map(lamdaA => P(9)(944),lamdaB => P(9)(946),s => s(9)(472),lamdaOut => P(8)(946));
U_G9947: entity G port map(lamdaA => P(9)(945),lamdaB => P(9)(947),s => s(9)(473),lamdaOut => P(8)(947));
U_F9948: entity F port map(lamdaA => P(9)(948),lamdaB => P(9)(950),lamdaOut => P(8)(948));
U_F9949: entity F port map(lamdaA => P(9)(949),lamdaB => P(9)(951),lamdaOut => P(8)(949));
U_G9950: entity G port map(lamdaA => P(9)(948),lamdaB => P(9)(950),s => s(9)(474),lamdaOut => P(8)(950));
U_G9951: entity G port map(lamdaA => P(9)(949),lamdaB => P(9)(951),s => s(9)(475),lamdaOut => P(8)(951));
U_F9952: entity F port map(lamdaA => P(9)(952),lamdaB => P(9)(954),lamdaOut => P(8)(952));
U_F9953: entity F port map(lamdaA => P(9)(953),lamdaB => P(9)(955),lamdaOut => P(8)(953));
U_G9954: entity G port map(lamdaA => P(9)(952),lamdaB => P(9)(954),s => s(9)(476),lamdaOut => P(8)(954));
U_G9955: entity G port map(lamdaA => P(9)(953),lamdaB => P(9)(955),s => s(9)(477),lamdaOut => P(8)(955));
U_F9956: entity F port map(lamdaA => P(9)(956),lamdaB => P(9)(958),lamdaOut => P(8)(956));
U_F9957: entity F port map(lamdaA => P(9)(957),lamdaB => P(9)(959),lamdaOut => P(8)(957));
U_G9958: entity G port map(lamdaA => P(9)(956),lamdaB => P(9)(958),s => s(9)(478),lamdaOut => P(8)(958));
U_G9959: entity G port map(lamdaA => P(9)(957),lamdaB => P(9)(959),s => s(9)(479),lamdaOut => P(8)(959));
U_F9960: entity F port map(lamdaA => P(9)(960),lamdaB => P(9)(962),lamdaOut => P(8)(960));
U_F9961: entity F port map(lamdaA => P(9)(961),lamdaB => P(9)(963),lamdaOut => P(8)(961));
U_G9962: entity G port map(lamdaA => P(9)(960),lamdaB => P(9)(962),s => s(9)(480),lamdaOut => P(8)(962));
U_G9963: entity G port map(lamdaA => P(9)(961),lamdaB => P(9)(963),s => s(9)(481),lamdaOut => P(8)(963));
U_F9964: entity F port map(lamdaA => P(9)(964),lamdaB => P(9)(966),lamdaOut => P(8)(964));
U_F9965: entity F port map(lamdaA => P(9)(965),lamdaB => P(9)(967),lamdaOut => P(8)(965));
U_G9966: entity G port map(lamdaA => P(9)(964),lamdaB => P(9)(966),s => s(9)(482),lamdaOut => P(8)(966));
U_G9967: entity G port map(lamdaA => P(9)(965),lamdaB => P(9)(967),s => s(9)(483),lamdaOut => P(8)(967));
U_F9968: entity F port map(lamdaA => P(9)(968),lamdaB => P(9)(970),lamdaOut => P(8)(968));
U_F9969: entity F port map(lamdaA => P(9)(969),lamdaB => P(9)(971),lamdaOut => P(8)(969));
U_G9970: entity G port map(lamdaA => P(9)(968),lamdaB => P(9)(970),s => s(9)(484),lamdaOut => P(8)(970));
U_G9971: entity G port map(lamdaA => P(9)(969),lamdaB => P(9)(971),s => s(9)(485),lamdaOut => P(8)(971));
U_F9972: entity F port map(lamdaA => P(9)(972),lamdaB => P(9)(974),lamdaOut => P(8)(972));
U_F9973: entity F port map(lamdaA => P(9)(973),lamdaB => P(9)(975),lamdaOut => P(8)(973));
U_G9974: entity G port map(lamdaA => P(9)(972),lamdaB => P(9)(974),s => s(9)(486),lamdaOut => P(8)(974));
U_G9975: entity G port map(lamdaA => P(9)(973),lamdaB => P(9)(975),s => s(9)(487),lamdaOut => P(8)(975));
U_F9976: entity F port map(lamdaA => P(9)(976),lamdaB => P(9)(978),lamdaOut => P(8)(976));
U_F9977: entity F port map(lamdaA => P(9)(977),lamdaB => P(9)(979),lamdaOut => P(8)(977));
U_G9978: entity G port map(lamdaA => P(9)(976),lamdaB => P(9)(978),s => s(9)(488),lamdaOut => P(8)(978));
U_G9979: entity G port map(lamdaA => P(9)(977),lamdaB => P(9)(979),s => s(9)(489),lamdaOut => P(8)(979));
U_F9980: entity F port map(lamdaA => P(9)(980),lamdaB => P(9)(982),lamdaOut => P(8)(980));
U_F9981: entity F port map(lamdaA => P(9)(981),lamdaB => P(9)(983),lamdaOut => P(8)(981));
U_G9982: entity G port map(lamdaA => P(9)(980),lamdaB => P(9)(982),s => s(9)(490),lamdaOut => P(8)(982));
U_G9983: entity G port map(lamdaA => P(9)(981),lamdaB => P(9)(983),s => s(9)(491),lamdaOut => P(8)(983));
U_F9984: entity F port map(lamdaA => P(9)(984),lamdaB => P(9)(986),lamdaOut => P(8)(984));
U_F9985: entity F port map(lamdaA => P(9)(985),lamdaB => P(9)(987),lamdaOut => P(8)(985));
U_G9986: entity G port map(lamdaA => P(9)(984),lamdaB => P(9)(986),s => s(9)(492),lamdaOut => P(8)(986));
U_G9987: entity G port map(lamdaA => P(9)(985),lamdaB => P(9)(987),s => s(9)(493),lamdaOut => P(8)(987));
U_F9988: entity F port map(lamdaA => P(9)(988),lamdaB => P(9)(990),lamdaOut => P(8)(988));
U_F9989: entity F port map(lamdaA => P(9)(989),lamdaB => P(9)(991),lamdaOut => P(8)(989));
U_G9990: entity G port map(lamdaA => P(9)(988),lamdaB => P(9)(990),s => s(9)(494),lamdaOut => P(8)(990));
U_G9991: entity G port map(lamdaA => P(9)(989),lamdaB => P(9)(991),s => s(9)(495),lamdaOut => P(8)(991));
U_F9992: entity F port map(lamdaA => P(9)(992),lamdaB => P(9)(994),lamdaOut => P(8)(992));
U_F9993: entity F port map(lamdaA => P(9)(993),lamdaB => P(9)(995),lamdaOut => P(8)(993));
U_G9994: entity G port map(lamdaA => P(9)(992),lamdaB => P(9)(994),s => s(9)(496),lamdaOut => P(8)(994));
U_G9995: entity G port map(lamdaA => P(9)(993),lamdaB => P(9)(995),s => s(9)(497),lamdaOut => P(8)(995));
U_F9996: entity F port map(lamdaA => P(9)(996),lamdaB => P(9)(998),lamdaOut => P(8)(996));
U_F9997: entity F port map(lamdaA => P(9)(997),lamdaB => P(9)(999),lamdaOut => P(8)(997));
U_G9998: entity G port map(lamdaA => P(9)(996),lamdaB => P(9)(998),s => s(9)(498),lamdaOut => P(8)(998));
U_G9999: entity G port map(lamdaA => P(9)(997),lamdaB => P(9)(999),s => s(9)(499),lamdaOut => P(8)(999));
U_F91000: entity F port map(lamdaA => P(9)(1000),lamdaB => P(9)(1002),lamdaOut => P(8)(1000));
U_F91001: entity F port map(lamdaA => P(9)(1001),lamdaB => P(9)(1003),lamdaOut => P(8)(1001));
U_G91002: entity G port map(lamdaA => P(9)(1000),lamdaB => P(9)(1002),s => s(9)(500),lamdaOut => P(8)(1002));
U_G91003: entity G port map(lamdaA => P(9)(1001),lamdaB => P(9)(1003),s => s(9)(501),lamdaOut => P(8)(1003));
U_F91004: entity F port map(lamdaA => P(9)(1004),lamdaB => P(9)(1006),lamdaOut => P(8)(1004));
U_F91005: entity F port map(lamdaA => P(9)(1005),lamdaB => P(9)(1007),lamdaOut => P(8)(1005));
U_G91006: entity G port map(lamdaA => P(9)(1004),lamdaB => P(9)(1006),s => s(9)(502),lamdaOut => P(8)(1006));
U_G91007: entity G port map(lamdaA => P(9)(1005),lamdaB => P(9)(1007),s => s(9)(503),lamdaOut => P(8)(1007));
U_F91008: entity F port map(lamdaA => P(9)(1008),lamdaB => P(9)(1010),lamdaOut => P(8)(1008));
U_F91009: entity F port map(lamdaA => P(9)(1009),lamdaB => P(9)(1011),lamdaOut => P(8)(1009));
U_G91010: entity G port map(lamdaA => P(9)(1008),lamdaB => P(9)(1010),s => s(9)(504),lamdaOut => P(8)(1010));
U_G91011: entity G port map(lamdaA => P(9)(1009),lamdaB => P(9)(1011),s => s(9)(505),lamdaOut => P(8)(1011));
U_F91012: entity F port map(lamdaA => P(9)(1012),lamdaB => P(9)(1014),lamdaOut => P(8)(1012));
U_F91013: entity F port map(lamdaA => P(9)(1013),lamdaB => P(9)(1015),lamdaOut => P(8)(1013));
U_G91014: entity G port map(lamdaA => P(9)(1012),lamdaB => P(9)(1014),s => s(9)(506),lamdaOut => P(8)(1014));
U_G91015: entity G port map(lamdaA => P(9)(1013),lamdaB => P(9)(1015),s => s(9)(507),lamdaOut => P(8)(1015));
U_F91016: entity F port map(lamdaA => P(9)(1016),lamdaB => P(9)(1018),lamdaOut => P(8)(1016));
U_F91017: entity F port map(lamdaA => P(9)(1017),lamdaB => P(9)(1019),lamdaOut => P(8)(1017));
U_G91018: entity G port map(lamdaA => P(9)(1016),lamdaB => P(9)(1018),s => s(9)(508),lamdaOut => P(8)(1018));
U_G91019: entity G port map(lamdaA => P(9)(1017),lamdaB => P(9)(1019),s => s(9)(509),lamdaOut => P(8)(1019));
U_F91020: entity F port map(lamdaA => P(9)(1020),lamdaB => P(9)(1022),lamdaOut => P(8)(1020));
U_F91021: entity F port map(lamdaA => P(9)(1021),lamdaB => P(9)(1023),lamdaOut => P(8)(1021));
U_G91022: entity G port map(lamdaA => P(9)(1020),lamdaB => P(9)(1022),s => s(9)(510),lamdaOut => P(8)(1022));
U_G91023: entity G port map(lamdaA => P(9)(1021),lamdaB => P(9)(1023),s => s(9)(511),lamdaOut => P(8)(1023));
-- STAGE 7
U_F80: entity F port map(lamdaA => P(8)(0),lamdaB => P(8)(4),lamdaOut => P(7)(0));
U_F81: entity F port map(lamdaA => P(8)(1),lamdaB => P(8)(5),lamdaOut => P(7)(1));
U_F82: entity F port map(lamdaA => P(8)(2),lamdaB => P(8)(6),lamdaOut => P(7)(2));
U_F83: entity F port map(lamdaA => P(8)(3),lamdaB => P(8)(7),lamdaOut => P(7)(3));
U_G84: entity G port map(lamdaA => P(8)(0),lamdaB => P(8)(4),s => s(8)(0),lamdaOut => P(7)(4));
U_G85: entity G port map(lamdaA => P(8)(1),lamdaB => P(8)(5),s => s(8)(1),lamdaOut => P(7)(5));
U_G86: entity G port map(lamdaA => P(8)(2),lamdaB => P(8)(6),s => s(8)(2),lamdaOut => P(7)(6));
U_G87: entity G port map(lamdaA => P(8)(3),lamdaB => P(8)(7),s => s(8)(3),lamdaOut => P(7)(7));
U_F88: entity F port map(lamdaA => P(8)(8),lamdaB => P(8)(12),lamdaOut => P(7)(8));
U_F89: entity F port map(lamdaA => P(8)(9),lamdaB => P(8)(13),lamdaOut => P(7)(9));
U_F810: entity F port map(lamdaA => P(8)(10),lamdaB => P(8)(14),lamdaOut => P(7)(10));
U_F811: entity F port map(lamdaA => P(8)(11),lamdaB => P(8)(15),lamdaOut => P(7)(11));
U_G812: entity G port map(lamdaA => P(8)(8),lamdaB => P(8)(12),s => s(8)(4),lamdaOut => P(7)(12));
U_G813: entity G port map(lamdaA => P(8)(9),lamdaB => P(8)(13),s => s(8)(5),lamdaOut => P(7)(13));
U_G814: entity G port map(lamdaA => P(8)(10),lamdaB => P(8)(14),s => s(8)(6),lamdaOut => P(7)(14));
U_G815: entity G port map(lamdaA => P(8)(11),lamdaB => P(8)(15),s => s(8)(7),lamdaOut => P(7)(15));
U_F816: entity F port map(lamdaA => P(8)(16),lamdaB => P(8)(20),lamdaOut => P(7)(16));
U_F817: entity F port map(lamdaA => P(8)(17),lamdaB => P(8)(21),lamdaOut => P(7)(17));
U_F818: entity F port map(lamdaA => P(8)(18),lamdaB => P(8)(22),lamdaOut => P(7)(18));
U_F819: entity F port map(lamdaA => P(8)(19),lamdaB => P(8)(23),lamdaOut => P(7)(19));
U_G820: entity G port map(lamdaA => P(8)(16),lamdaB => P(8)(20),s => s(8)(8),lamdaOut => P(7)(20));
U_G821: entity G port map(lamdaA => P(8)(17),lamdaB => P(8)(21),s => s(8)(9),lamdaOut => P(7)(21));
U_G822: entity G port map(lamdaA => P(8)(18),lamdaB => P(8)(22),s => s(8)(10),lamdaOut => P(7)(22));
U_G823: entity G port map(lamdaA => P(8)(19),lamdaB => P(8)(23),s => s(8)(11),lamdaOut => P(7)(23));
U_F824: entity F port map(lamdaA => P(8)(24),lamdaB => P(8)(28),lamdaOut => P(7)(24));
U_F825: entity F port map(lamdaA => P(8)(25),lamdaB => P(8)(29),lamdaOut => P(7)(25));
U_F826: entity F port map(lamdaA => P(8)(26),lamdaB => P(8)(30),lamdaOut => P(7)(26));
U_F827: entity F port map(lamdaA => P(8)(27),lamdaB => P(8)(31),lamdaOut => P(7)(27));
U_G828: entity G port map(lamdaA => P(8)(24),lamdaB => P(8)(28),s => s(8)(12),lamdaOut => P(7)(28));
U_G829: entity G port map(lamdaA => P(8)(25),lamdaB => P(8)(29),s => s(8)(13),lamdaOut => P(7)(29));
U_G830: entity G port map(lamdaA => P(8)(26),lamdaB => P(8)(30),s => s(8)(14),lamdaOut => P(7)(30));
U_G831: entity G port map(lamdaA => P(8)(27),lamdaB => P(8)(31),s => s(8)(15),lamdaOut => P(7)(31));
U_F832: entity F port map(lamdaA => P(8)(32),lamdaB => P(8)(36),lamdaOut => P(7)(32));
U_F833: entity F port map(lamdaA => P(8)(33),lamdaB => P(8)(37),lamdaOut => P(7)(33));
U_F834: entity F port map(lamdaA => P(8)(34),lamdaB => P(8)(38),lamdaOut => P(7)(34));
U_F835: entity F port map(lamdaA => P(8)(35),lamdaB => P(8)(39),lamdaOut => P(7)(35));
U_G836: entity G port map(lamdaA => P(8)(32),lamdaB => P(8)(36),s => s(8)(16),lamdaOut => P(7)(36));
U_G837: entity G port map(lamdaA => P(8)(33),lamdaB => P(8)(37),s => s(8)(17),lamdaOut => P(7)(37));
U_G838: entity G port map(lamdaA => P(8)(34),lamdaB => P(8)(38),s => s(8)(18),lamdaOut => P(7)(38));
U_G839: entity G port map(lamdaA => P(8)(35),lamdaB => P(8)(39),s => s(8)(19),lamdaOut => P(7)(39));
U_F840: entity F port map(lamdaA => P(8)(40),lamdaB => P(8)(44),lamdaOut => P(7)(40));
U_F841: entity F port map(lamdaA => P(8)(41),lamdaB => P(8)(45),lamdaOut => P(7)(41));
U_F842: entity F port map(lamdaA => P(8)(42),lamdaB => P(8)(46),lamdaOut => P(7)(42));
U_F843: entity F port map(lamdaA => P(8)(43),lamdaB => P(8)(47),lamdaOut => P(7)(43));
U_G844: entity G port map(lamdaA => P(8)(40),lamdaB => P(8)(44),s => s(8)(20),lamdaOut => P(7)(44));
U_G845: entity G port map(lamdaA => P(8)(41),lamdaB => P(8)(45),s => s(8)(21),lamdaOut => P(7)(45));
U_G846: entity G port map(lamdaA => P(8)(42),lamdaB => P(8)(46),s => s(8)(22),lamdaOut => P(7)(46));
U_G847: entity G port map(lamdaA => P(8)(43),lamdaB => P(8)(47),s => s(8)(23),lamdaOut => P(7)(47));
U_F848: entity F port map(lamdaA => P(8)(48),lamdaB => P(8)(52),lamdaOut => P(7)(48));
U_F849: entity F port map(lamdaA => P(8)(49),lamdaB => P(8)(53),lamdaOut => P(7)(49));
U_F850: entity F port map(lamdaA => P(8)(50),lamdaB => P(8)(54),lamdaOut => P(7)(50));
U_F851: entity F port map(lamdaA => P(8)(51),lamdaB => P(8)(55),lamdaOut => P(7)(51));
U_G852: entity G port map(lamdaA => P(8)(48),lamdaB => P(8)(52),s => s(8)(24),lamdaOut => P(7)(52));
U_G853: entity G port map(lamdaA => P(8)(49),lamdaB => P(8)(53),s => s(8)(25),lamdaOut => P(7)(53));
U_G854: entity G port map(lamdaA => P(8)(50),lamdaB => P(8)(54),s => s(8)(26),lamdaOut => P(7)(54));
U_G855: entity G port map(lamdaA => P(8)(51),lamdaB => P(8)(55),s => s(8)(27),lamdaOut => P(7)(55));
U_F856: entity F port map(lamdaA => P(8)(56),lamdaB => P(8)(60),lamdaOut => P(7)(56));
U_F857: entity F port map(lamdaA => P(8)(57),lamdaB => P(8)(61),lamdaOut => P(7)(57));
U_F858: entity F port map(lamdaA => P(8)(58),lamdaB => P(8)(62),lamdaOut => P(7)(58));
U_F859: entity F port map(lamdaA => P(8)(59),lamdaB => P(8)(63),lamdaOut => P(7)(59));
U_G860: entity G port map(lamdaA => P(8)(56),lamdaB => P(8)(60),s => s(8)(28),lamdaOut => P(7)(60));
U_G861: entity G port map(lamdaA => P(8)(57),lamdaB => P(8)(61),s => s(8)(29),lamdaOut => P(7)(61));
U_G862: entity G port map(lamdaA => P(8)(58),lamdaB => P(8)(62),s => s(8)(30),lamdaOut => P(7)(62));
U_G863: entity G port map(lamdaA => P(8)(59),lamdaB => P(8)(63),s => s(8)(31),lamdaOut => P(7)(63));
U_F864: entity F port map(lamdaA => P(8)(64),lamdaB => P(8)(68),lamdaOut => P(7)(64));
U_F865: entity F port map(lamdaA => P(8)(65),lamdaB => P(8)(69),lamdaOut => P(7)(65));
U_F866: entity F port map(lamdaA => P(8)(66),lamdaB => P(8)(70),lamdaOut => P(7)(66));
U_F867: entity F port map(lamdaA => P(8)(67),lamdaB => P(8)(71),lamdaOut => P(7)(67));
U_G868: entity G port map(lamdaA => P(8)(64),lamdaB => P(8)(68),s => s(8)(32),lamdaOut => P(7)(68));
U_G869: entity G port map(lamdaA => P(8)(65),lamdaB => P(8)(69),s => s(8)(33),lamdaOut => P(7)(69));
U_G870: entity G port map(lamdaA => P(8)(66),lamdaB => P(8)(70),s => s(8)(34),lamdaOut => P(7)(70));
U_G871: entity G port map(lamdaA => P(8)(67),lamdaB => P(8)(71),s => s(8)(35),lamdaOut => P(7)(71));
U_F872: entity F port map(lamdaA => P(8)(72),lamdaB => P(8)(76),lamdaOut => P(7)(72));
U_F873: entity F port map(lamdaA => P(8)(73),lamdaB => P(8)(77),lamdaOut => P(7)(73));
U_F874: entity F port map(lamdaA => P(8)(74),lamdaB => P(8)(78),lamdaOut => P(7)(74));
U_F875: entity F port map(lamdaA => P(8)(75),lamdaB => P(8)(79),lamdaOut => P(7)(75));
U_G876: entity G port map(lamdaA => P(8)(72),lamdaB => P(8)(76),s => s(8)(36),lamdaOut => P(7)(76));
U_G877: entity G port map(lamdaA => P(8)(73),lamdaB => P(8)(77),s => s(8)(37),lamdaOut => P(7)(77));
U_G878: entity G port map(lamdaA => P(8)(74),lamdaB => P(8)(78),s => s(8)(38),lamdaOut => P(7)(78));
U_G879: entity G port map(lamdaA => P(8)(75),lamdaB => P(8)(79),s => s(8)(39),lamdaOut => P(7)(79));
U_F880: entity F port map(lamdaA => P(8)(80),lamdaB => P(8)(84),lamdaOut => P(7)(80));
U_F881: entity F port map(lamdaA => P(8)(81),lamdaB => P(8)(85),lamdaOut => P(7)(81));
U_F882: entity F port map(lamdaA => P(8)(82),lamdaB => P(8)(86),lamdaOut => P(7)(82));
U_F883: entity F port map(lamdaA => P(8)(83),lamdaB => P(8)(87),lamdaOut => P(7)(83));
U_G884: entity G port map(lamdaA => P(8)(80),lamdaB => P(8)(84),s => s(8)(40),lamdaOut => P(7)(84));
U_G885: entity G port map(lamdaA => P(8)(81),lamdaB => P(8)(85),s => s(8)(41),lamdaOut => P(7)(85));
U_G886: entity G port map(lamdaA => P(8)(82),lamdaB => P(8)(86),s => s(8)(42),lamdaOut => P(7)(86));
U_G887: entity G port map(lamdaA => P(8)(83),lamdaB => P(8)(87),s => s(8)(43),lamdaOut => P(7)(87));
U_F888: entity F port map(lamdaA => P(8)(88),lamdaB => P(8)(92),lamdaOut => P(7)(88));
U_F889: entity F port map(lamdaA => P(8)(89),lamdaB => P(8)(93),lamdaOut => P(7)(89));
U_F890: entity F port map(lamdaA => P(8)(90),lamdaB => P(8)(94),lamdaOut => P(7)(90));
U_F891: entity F port map(lamdaA => P(8)(91),lamdaB => P(8)(95),lamdaOut => P(7)(91));
U_G892: entity G port map(lamdaA => P(8)(88),lamdaB => P(8)(92),s => s(8)(44),lamdaOut => P(7)(92));
U_G893: entity G port map(lamdaA => P(8)(89),lamdaB => P(8)(93),s => s(8)(45),lamdaOut => P(7)(93));
U_G894: entity G port map(lamdaA => P(8)(90),lamdaB => P(8)(94),s => s(8)(46),lamdaOut => P(7)(94));
U_G895: entity G port map(lamdaA => P(8)(91),lamdaB => P(8)(95),s => s(8)(47),lamdaOut => P(7)(95));
U_F896: entity F port map(lamdaA => P(8)(96),lamdaB => P(8)(100),lamdaOut => P(7)(96));
U_F897: entity F port map(lamdaA => P(8)(97),lamdaB => P(8)(101),lamdaOut => P(7)(97));
U_F898: entity F port map(lamdaA => P(8)(98),lamdaB => P(8)(102),lamdaOut => P(7)(98));
U_F899: entity F port map(lamdaA => P(8)(99),lamdaB => P(8)(103),lamdaOut => P(7)(99));
U_G8100: entity G port map(lamdaA => P(8)(96),lamdaB => P(8)(100),s => s(8)(48),lamdaOut => P(7)(100));
U_G8101: entity G port map(lamdaA => P(8)(97),lamdaB => P(8)(101),s => s(8)(49),lamdaOut => P(7)(101));
U_G8102: entity G port map(lamdaA => P(8)(98),lamdaB => P(8)(102),s => s(8)(50),lamdaOut => P(7)(102));
U_G8103: entity G port map(lamdaA => P(8)(99),lamdaB => P(8)(103),s => s(8)(51),lamdaOut => P(7)(103));
U_F8104: entity F port map(lamdaA => P(8)(104),lamdaB => P(8)(108),lamdaOut => P(7)(104));
U_F8105: entity F port map(lamdaA => P(8)(105),lamdaB => P(8)(109),lamdaOut => P(7)(105));
U_F8106: entity F port map(lamdaA => P(8)(106),lamdaB => P(8)(110),lamdaOut => P(7)(106));
U_F8107: entity F port map(lamdaA => P(8)(107),lamdaB => P(8)(111),lamdaOut => P(7)(107));
U_G8108: entity G port map(lamdaA => P(8)(104),lamdaB => P(8)(108),s => s(8)(52),lamdaOut => P(7)(108));
U_G8109: entity G port map(lamdaA => P(8)(105),lamdaB => P(8)(109),s => s(8)(53),lamdaOut => P(7)(109));
U_G8110: entity G port map(lamdaA => P(8)(106),lamdaB => P(8)(110),s => s(8)(54),lamdaOut => P(7)(110));
U_G8111: entity G port map(lamdaA => P(8)(107),lamdaB => P(8)(111),s => s(8)(55),lamdaOut => P(7)(111));
U_F8112: entity F port map(lamdaA => P(8)(112),lamdaB => P(8)(116),lamdaOut => P(7)(112));
U_F8113: entity F port map(lamdaA => P(8)(113),lamdaB => P(8)(117),lamdaOut => P(7)(113));
U_F8114: entity F port map(lamdaA => P(8)(114),lamdaB => P(8)(118),lamdaOut => P(7)(114));
U_F8115: entity F port map(lamdaA => P(8)(115),lamdaB => P(8)(119),lamdaOut => P(7)(115));
U_G8116: entity G port map(lamdaA => P(8)(112),lamdaB => P(8)(116),s => s(8)(56),lamdaOut => P(7)(116));
U_G8117: entity G port map(lamdaA => P(8)(113),lamdaB => P(8)(117),s => s(8)(57),lamdaOut => P(7)(117));
U_G8118: entity G port map(lamdaA => P(8)(114),lamdaB => P(8)(118),s => s(8)(58),lamdaOut => P(7)(118));
U_G8119: entity G port map(lamdaA => P(8)(115),lamdaB => P(8)(119),s => s(8)(59),lamdaOut => P(7)(119));
U_F8120: entity F port map(lamdaA => P(8)(120),lamdaB => P(8)(124),lamdaOut => P(7)(120));
U_F8121: entity F port map(lamdaA => P(8)(121),lamdaB => P(8)(125),lamdaOut => P(7)(121));
U_F8122: entity F port map(lamdaA => P(8)(122),lamdaB => P(8)(126),lamdaOut => P(7)(122));
U_F8123: entity F port map(lamdaA => P(8)(123),lamdaB => P(8)(127),lamdaOut => P(7)(123));
U_G8124: entity G port map(lamdaA => P(8)(120),lamdaB => P(8)(124),s => s(8)(60),lamdaOut => P(7)(124));
U_G8125: entity G port map(lamdaA => P(8)(121),lamdaB => P(8)(125),s => s(8)(61),lamdaOut => P(7)(125));
U_G8126: entity G port map(lamdaA => P(8)(122),lamdaB => P(8)(126),s => s(8)(62),lamdaOut => P(7)(126));
U_G8127: entity G port map(lamdaA => P(8)(123),lamdaB => P(8)(127),s => s(8)(63),lamdaOut => P(7)(127));
U_F8128: entity F port map(lamdaA => P(8)(128),lamdaB => P(8)(132),lamdaOut => P(7)(128));
U_F8129: entity F port map(lamdaA => P(8)(129),lamdaB => P(8)(133),lamdaOut => P(7)(129));
U_F8130: entity F port map(lamdaA => P(8)(130),lamdaB => P(8)(134),lamdaOut => P(7)(130));
U_F8131: entity F port map(lamdaA => P(8)(131),lamdaB => P(8)(135),lamdaOut => P(7)(131));
U_G8132: entity G port map(lamdaA => P(8)(128),lamdaB => P(8)(132),s => s(8)(64),lamdaOut => P(7)(132));
U_G8133: entity G port map(lamdaA => P(8)(129),lamdaB => P(8)(133),s => s(8)(65),lamdaOut => P(7)(133));
U_G8134: entity G port map(lamdaA => P(8)(130),lamdaB => P(8)(134),s => s(8)(66),lamdaOut => P(7)(134));
U_G8135: entity G port map(lamdaA => P(8)(131),lamdaB => P(8)(135),s => s(8)(67),lamdaOut => P(7)(135));
U_F8136: entity F port map(lamdaA => P(8)(136),lamdaB => P(8)(140),lamdaOut => P(7)(136));
U_F8137: entity F port map(lamdaA => P(8)(137),lamdaB => P(8)(141),lamdaOut => P(7)(137));
U_F8138: entity F port map(lamdaA => P(8)(138),lamdaB => P(8)(142),lamdaOut => P(7)(138));
U_F8139: entity F port map(lamdaA => P(8)(139),lamdaB => P(8)(143),lamdaOut => P(7)(139));
U_G8140: entity G port map(lamdaA => P(8)(136),lamdaB => P(8)(140),s => s(8)(68),lamdaOut => P(7)(140));
U_G8141: entity G port map(lamdaA => P(8)(137),lamdaB => P(8)(141),s => s(8)(69),lamdaOut => P(7)(141));
U_G8142: entity G port map(lamdaA => P(8)(138),lamdaB => P(8)(142),s => s(8)(70),lamdaOut => P(7)(142));
U_G8143: entity G port map(lamdaA => P(8)(139),lamdaB => P(8)(143),s => s(8)(71),lamdaOut => P(7)(143));
U_F8144: entity F port map(lamdaA => P(8)(144),lamdaB => P(8)(148),lamdaOut => P(7)(144));
U_F8145: entity F port map(lamdaA => P(8)(145),lamdaB => P(8)(149),lamdaOut => P(7)(145));
U_F8146: entity F port map(lamdaA => P(8)(146),lamdaB => P(8)(150),lamdaOut => P(7)(146));
U_F8147: entity F port map(lamdaA => P(8)(147),lamdaB => P(8)(151),lamdaOut => P(7)(147));
U_G8148: entity G port map(lamdaA => P(8)(144),lamdaB => P(8)(148),s => s(8)(72),lamdaOut => P(7)(148));
U_G8149: entity G port map(lamdaA => P(8)(145),lamdaB => P(8)(149),s => s(8)(73),lamdaOut => P(7)(149));
U_G8150: entity G port map(lamdaA => P(8)(146),lamdaB => P(8)(150),s => s(8)(74),lamdaOut => P(7)(150));
U_G8151: entity G port map(lamdaA => P(8)(147),lamdaB => P(8)(151),s => s(8)(75),lamdaOut => P(7)(151));
U_F8152: entity F port map(lamdaA => P(8)(152),lamdaB => P(8)(156),lamdaOut => P(7)(152));
U_F8153: entity F port map(lamdaA => P(8)(153),lamdaB => P(8)(157),lamdaOut => P(7)(153));
U_F8154: entity F port map(lamdaA => P(8)(154),lamdaB => P(8)(158),lamdaOut => P(7)(154));
U_F8155: entity F port map(lamdaA => P(8)(155),lamdaB => P(8)(159),lamdaOut => P(7)(155));
U_G8156: entity G port map(lamdaA => P(8)(152),lamdaB => P(8)(156),s => s(8)(76),lamdaOut => P(7)(156));
U_G8157: entity G port map(lamdaA => P(8)(153),lamdaB => P(8)(157),s => s(8)(77),lamdaOut => P(7)(157));
U_G8158: entity G port map(lamdaA => P(8)(154),lamdaB => P(8)(158),s => s(8)(78),lamdaOut => P(7)(158));
U_G8159: entity G port map(lamdaA => P(8)(155),lamdaB => P(8)(159),s => s(8)(79),lamdaOut => P(7)(159));
U_F8160: entity F port map(lamdaA => P(8)(160),lamdaB => P(8)(164),lamdaOut => P(7)(160));
U_F8161: entity F port map(lamdaA => P(8)(161),lamdaB => P(8)(165),lamdaOut => P(7)(161));
U_F8162: entity F port map(lamdaA => P(8)(162),lamdaB => P(8)(166),lamdaOut => P(7)(162));
U_F8163: entity F port map(lamdaA => P(8)(163),lamdaB => P(8)(167),lamdaOut => P(7)(163));
U_G8164: entity G port map(lamdaA => P(8)(160),lamdaB => P(8)(164),s => s(8)(80),lamdaOut => P(7)(164));
U_G8165: entity G port map(lamdaA => P(8)(161),lamdaB => P(8)(165),s => s(8)(81),lamdaOut => P(7)(165));
U_G8166: entity G port map(lamdaA => P(8)(162),lamdaB => P(8)(166),s => s(8)(82),lamdaOut => P(7)(166));
U_G8167: entity G port map(lamdaA => P(8)(163),lamdaB => P(8)(167),s => s(8)(83),lamdaOut => P(7)(167));
U_F8168: entity F port map(lamdaA => P(8)(168),lamdaB => P(8)(172),lamdaOut => P(7)(168));
U_F8169: entity F port map(lamdaA => P(8)(169),lamdaB => P(8)(173),lamdaOut => P(7)(169));
U_F8170: entity F port map(lamdaA => P(8)(170),lamdaB => P(8)(174),lamdaOut => P(7)(170));
U_F8171: entity F port map(lamdaA => P(8)(171),lamdaB => P(8)(175),lamdaOut => P(7)(171));
U_G8172: entity G port map(lamdaA => P(8)(168),lamdaB => P(8)(172),s => s(8)(84),lamdaOut => P(7)(172));
U_G8173: entity G port map(lamdaA => P(8)(169),lamdaB => P(8)(173),s => s(8)(85),lamdaOut => P(7)(173));
U_G8174: entity G port map(lamdaA => P(8)(170),lamdaB => P(8)(174),s => s(8)(86),lamdaOut => P(7)(174));
U_G8175: entity G port map(lamdaA => P(8)(171),lamdaB => P(8)(175),s => s(8)(87),lamdaOut => P(7)(175));
U_F8176: entity F port map(lamdaA => P(8)(176),lamdaB => P(8)(180),lamdaOut => P(7)(176));
U_F8177: entity F port map(lamdaA => P(8)(177),lamdaB => P(8)(181),lamdaOut => P(7)(177));
U_F8178: entity F port map(lamdaA => P(8)(178),lamdaB => P(8)(182),lamdaOut => P(7)(178));
U_F8179: entity F port map(lamdaA => P(8)(179),lamdaB => P(8)(183),lamdaOut => P(7)(179));
U_G8180: entity G port map(lamdaA => P(8)(176),lamdaB => P(8)(180),s => s(8)(88),lamdaOut => P(7)(180));
U_G8181: entity G port map(lamdaA => P(8)(177),lamdaB => P(8)(181),s => s(8)(89),lamdaOut => P(7)(181));
U_G8182: entity G port map(lamdaA => P(8)(178),lamdaB => P(8)(182),s => s(8)(90),lamdaOut => P(7)(182));
U_G8183: entity G port map(lamdaA => P(8)(179),lamdaB => P(8)(183),s => s(8)(91),lamdaOut => P(7)(183));
U_F8184: entity F port map(lamdaA => P(8)(184),lamdaB => P(8)(188),lamdaOut => P(7)(184));
U_F8185: entity F port map(lamdaA => P(8)(185),lamdaB => P(8)(189),lamdaOut => P(7)(185));
U_F8186: entity F port map(lamdaA => P(8)(186),lamdaB => P(8)(190),lamdaOut => P(7)(186));
U_F8187: entity F port map(lamdaA => P(8)(187),lamdaB => P(8)(191),lamdaOut => P(7)(187));
U_G8188: entity G port map(lamdaA => P(8)(184),lamdaB => P(8)(188),s => s(8)(92),lamdaOut => P(7)(188));
U_G8189: entity G port map(lamdaA => P(8)(185),lamdaB => P(8)(189),s => s(8)(93),lamdaOut => P(7)(189));
U_G8190: entity G port map(lamdaA => P(8)(186),lamdaB => P(8)(190),s => s(8)(94),lamdaOut => P(7)(190));
U_G8191: entity G port map(lamdaA => P(8)(187),lamdaB => P(8)(191),s => s(8)(95),lamdaOut => P(7)(191));
U_F8192: entity F port map(lamdaA => P(8)(192),lamdaB => P(8)(196),lamdaOut => P(7)(192));
U_F8193: entity F port map(lamdaA => P(8)(193),lamdaB => P(8)(197),lamdaOut => P(7)(193));
U_F8194: entity F port map(lamdaA => P(8)(194),lamdaB => P(8)(198),lamdaOut => P(7)(194));
U_F8195: entity F port map(lamdaA => P(8)(195),lamdaB => P(8)(199),lamdaOut => P(7)(195));
U_G8196: entity G port map(lamdaA => P(8)(192),lamdaB => P(8)(196),s => s(8)(96),lamdaOut => P(7)(196));
U_G8197: entity G port map(lamdaA => P(8)(193),lamdaB => P(8)(197),s => s(8)(97),lamdaOut => P(7)(197));
U_G8198: entity G port map(lamdaA => P(8)(194),lamdaB => P(8)(198),s => s(8)(98),lamdaOut => P(7)(198));
U_G8199: entity G port map(lamdaA => P(8)(195),lamdaB => P(8)(199),s => s(8)(99),lamdaOut => P(7)(199));
U_F8200: entity F port map(lamdaA => P(8)(200),lamdaB => P(8)(204),lamdaOut => P(7)(200));
U_F8201: entity F port map(lamdaA => P(8)(201),lamdaB => P(8)(205),lamdaOut => P(7)(201));
U_F8202: entity F port map(lamdaA => P(8)(202),lamdaB => P(8)(206),lamdaOut => P(7)(202));
U_F8203: entity F port map(lamdaA => P(8)(203),lamdaB => P(8)(207),lamdaOut => P(7)(203));
U_G8204: entity G port map(lamdaA => P(8)(200),lamdaB => P(8)(204),s => s(8)(100),lamdaOut => P(7)(204));
U_G8205: entity G port map(lamdaA => P(8)(201),lamdaB => P(8)(205),s => s(8)(101),lamdaOut => P(7)(205));
U_G8206: entity G port map(lamdaA => P(8)(202),lamdaB => P(8)(206),s => s(8)(102),lamdaOut => P(7)(206));
U_G8207: entity G port map(lamdaA => P(8)(203),lamdaB => P(8)(207),s => s(8)(103),lamdaOut => P(7)(207));
U_F8208: entity F port map(lamdaA => P(8)(208),lamdaB => P(8)(212),lamdaOut => P(7)(208));
U_F8209: entity F port map(lamdaA => P(8)(209),lamdaB => P(8)(213),lamdaOut => P(7)(209));
U_F8210: entity F port map(lamdaA => P(8)(210),lamdaB => P(8)(214),lamdaOut => P(7)(210));
U_F8211: entity F port map(lamdaA => P(8)(211),lamdaB => P(8)(215),lamdaOut => P(7)(211));
U_G8212: entity G port map(lamdaA => P(8)(208),lamdaB => P(8)(212),s => s(8)(104),lamdaOut => P(7)(212));
U_G8213: entity G port map(lamdaA => P(8)(209),lamdaB => P(8)(213),s => s(8)(105),lamdaOut => P(7)(213));
U_G8214: entity G port map(lamdaA => P(8)(210),lamdaB => P(8)(214),s => s(8)(106),lamdaOut => P(7)(214));
U_G8215: entity G port map(lamdaA => P(8)(211),lamdaB => P(8)(215),s => s(8)(107),lamdaOut => P(7)(215));
U_F8216: entity F port map(lamdaA => P(8)(216),lamdaB => P(8)(220),lamdaOut => P(7)(216));
U_F8217: entity F port map(lamdaA => P(8)(217),lamdaB => P(8)(221),lamdaOut => P(7)(217));
U_F8218: entity F port map(lamdaA => P(8)(218),lamdaB => P(8)(222),lamdaOut => P(7)(218));
U_F8219: entity F port map(lamdaA => P(8)(219),lamdaB => P(8)(223),lamdaOut => P(7)(219));
U_G8220: entity G port map(lamdaA => P(8)(216),lamdaB => P(8)(220),s => s(8)(108),lamdaOut => P(7)(220));
U_G8221: entity G port map(lamdaA => P(8)(217),lamdaB => P(8)(221),s => s(8)(109),lamdaOut => P(7)(221));
U_G8222: entity G port map(lamdaA => P(8)(218),lamdaB => P(8)(222),s => s(8)(110),lamdaOut => P(7)(222));
U_G8223: entity G port map(lamdaA => P(8)(219),lamdaB => P(8)(223),s => s(8)(111),lamdaOut => P(7)(223));
U_F8224: entity F port map(lamdaA => P(8)(224),lamdaB => P(8)(228),lamdaOut => P(7)(224));
U_F8225: entity F port map(lamdaA => P(8)(225),lamdaB => P(8)(229),lamdaOut => P(7)(225));
U_F8226: entity F port map(lamdaA => P(8)(226),lamdaB => P(8)(230),lamdaOut => P(7)(226));
U_F8227: entity F port map(lamdaA => P(8)(227),lamdaB => P(8)(231),lamdaOut => P(7)(227));
U_G8228: entity G port map(lamdaA => P(8)(224),lamdaB => P(8)(228),s => s(8)(112),lamdaOut => P(7)(228));
U_G8229: entity G port map(lamdaA => P(8)(225),lamdaB => P(8)(229),s => s(8)(113),lamdaOut => P(7)(229));
U_G8230: entity G port map(lamdaA => P(8)(226),lamdaB => P(8)(230),s => s(8)(114),lamdaOut => P(7)(230));
U_G8231: entity G port map(lamdaA => P(8)(227),lamdaB => P(8)(231),s => s(8)(115),lamdaOut => P(7)(231));
U_F8232: entity F port map(lamdaA => P(8)(232),lamdaB => P(8)(236),lamdaOut => P(7)(232));
U_F8233: entity F port map(lamdaA => P(8)(233),lamdaB => P(8)(237),lamdaOut => P(7)(233));
U_F8234: entity F port map(lamdaA => P(8)(234),lamdaB => P(8)(238),lamdaOut => P(7)(234));
U_F8235: entity F port map(lamdaA => P(8)(235),lamdaB => P(8)(239),lamdaOut => P(7)(235));
U_G8236: entity G port map(lamdaA => P(8)(232),lamdaB => P(8)(236),s => s(8)(116),lamdaOut => P(7)(236));
U_G8237: entity G port map(lamdaA => P(8)(233),lamdaB => P(8)(237),s => s(8)(117),lamdaOut => P(7)(237));
U_G8238: entity G port map(lamdaA => P(8)(234),lamdaB => P(8)(238),s => s(8)(118),lamdaOut => P(7)(238));
U_G8239: entity G port map(lamdaA => P(8)(235),lamdaB => P(8)(239),s => s(8)(119),lamdaOut => P(7)(239));
U_F8240: entity F port map(lamdaA => P(8)(240),lamdaB => P(8)(244),lamdaOut => P(7)(240));
U_F8241: entity F port map(lamdaA => P(8)(241),lamdaB => P(8)(245),lamdaOut => P(7)(241));
U_F8242: entity F port map(lamdaA => P(8)(242),lamdaB => P(8)(246),lamdaOut => P(7)(242));
U_F8243: entity F port map(lamdaA => P(8)(243),lamdaB => P(8)(247),lamdaOut => P(7)(243));
U_G8244: entity G port map(lamdaA => P(8)(240),lamdaB => P(8)(244),s => s(8)(120),lamdaOut => P(7)(244));
U_G8245: entity G port map(lamdaA => P(8)(241),lamdaB => P(8)(245),s => s(8)(121),lamdaOut => P(7)(245));
U_G8246: entity G port map(lamdaA => P(8)(242),lamdaB => P(8)(246),s => s(8)(122),lamdaOut => P(7)(246));
U_G8247: entity G port map(lamdaA => P(8)(243),lamdaB => P(8)(247),s => s(8)(123),lamdaOut => P(7)(247));
U_F8248: entity F port map(lamdaA => P(8)(248),lamdaB => P(8)(252),lamdaOut => P(7)(248));
U_F8249: entity F port map(lamdaA => P(8)(249),lamdaB => P(8)(253),lamdaOut => P(7)(249));
U_F8250: entity F port map(lamdaA => P(8)(250),lamdaB => P(8)(254),lamdaOut => P(7)(250));
U_F8251: entity F port map(lamdaA => P(8)(251),lamdaB => P(8)(255),lamdaOut => P(7)(251));
U_G8252: entity G port map(lamdaA => P(8)(248),lamdaB => P(8)(252),s => s(8)(124),lamdaOut => P(7)(252));
U_G8253: entity G port map(lamdaA => P(8)(249),lamdaB => P(8)(253),s => s(8)(125),lamdaOut => P(7)(253));
U_G8254: entity G port map(lamdaA => P(8)(250),lamdaB => P(8)(254),s => s(8)(126),lamdaOut => P(7)(254));
U_G8255: entity G port map(lamdaA => P(8)(251),lamdaB => P(8)(255),s => s(8)(127),lamdaOut => P(7)(255));
U_F8256: entity F port map(lamdaA => P(8)(256),lamdaB => P(8)(260),lamdaOut => P(7)(256));
U_F8257: entity F port map(lamdaA => P(8)(257),lamdaB => P(8)(261),lamdaOut => P(7)(257));
U_F8258: entity F port map(lamdaA => P(8)(258),lamdaB => P(8)(262),lamdaOut => P(7)(258));
U_F8259: entity F port map(lamdaA => P(8)(259),lamdaB => P(8)(263),lamdaOut => P(7)(259));
U_G8260: entity G port map(lamdaA => P(8)(256),lamdaB => P(8)(260),s => s(8)(128),lamdaOut => P(7)(260));
U_G8261: entity G port map(lamdaA => P(8)(257),lamdaB => P(8)(261),s => s(8)(129),lamdaOut => P(7)(261));
U_G8262: entity G port map(lamdaA => P(8)(258),lamdaB => P(8)(262),s => s(8)(130),lamdaOut => P(7)(262));
U_G8263: entity G port map(lamdaA => P(8)(259),lamdaB => P(8)(263),s => s(8)(131),lamdaOut => P(7)(263));
U_F8264: entity F port map(lamdaA => P(8)(264),lamdaB => P(8)(268),lamdaOut => P(7)(264));
U_F8265: entity F port map(lamdaA => P(8)(265),lamdaB => P(8)(269),lamdaOut => P(7)(265));
U_F8266: entity F port map(lamdaA => P(8)(266),lamdaB => P(8)(270),lamdaOut => P(7)(266));
U_F8267: entity F port map(lamdaA => P(8)(267),lamdaB => P(8)(271),lamdaOut => P(7)(267));
U_G8268: entity G port map(lamdaA => P(8)(264),lamdaB => P(8)(268),s => s(8)(132),lamdaOut => P(7)(268));
U_G8269: entity G port map(lamdaA => P(8)(265),lamdaB => P(8)(269),s => s(8)(133),lamdaOut => P(7)(269));
U_G8270: entity G port map(lamdaA => P(8)(266),lamdaB => P(8)(270),s => s(8)(134),lamdaOut => P(7)(270));
U_G8271: entity G port map(lamdaA => P(8)(267),lamdaB => P(8)(271),s => s(8)(135),lamdaOut => P(7)(271));
U_F8272: entity F port map(lamdaA => P(8)(272),lamdaB => P(8)(276),lamdaOut => P(7)(272));
U_F8273: entity F port map(lamdaA => P(8)(273),lamdaB => P(8)(277),lamdaOut => P(7)(273));
U_F8274: entity F port map(lamdaA => P(8)(274),lamdaB => P(8)(278),lamdaOut => P(7)(274));
U_F8275: entity F port map(lamdaA => P(8)(275),lamdaB => P(8)(279),lamdaOut => P(7)(275));
U_G8276: entity G port map(lamdaA => P(8)(272),lamdaB => P(8)(276),s => s(8)(136),lamdaOut => P(7)(276));
U_G8277: entity G port map(lamdaA => P(8)(273),lamdaB => P(8)(277),s => s(8)(137),lamdaOut => P(7)(277));
U_G8278: entity G port map(lamdaA => P(8)(274),lamdaB => P(8)(278),s => s(8)(138),lamdaOut => P(7)(278));
U_G8279: entity G port map(lamdaA => P(8)(275),lamdaB => P(8)(279),s => s(8)(139),lamdaOut => P(7)(279));
U_F8280: entity F port map(lamdaA => P(8)(280),lamdaB => P(8)(284),lamdaOut => P(7)(280));
U_F8281: entity F port map(lamdaA => P(8)(281),lamdaB => P(8)(285),lamdaOut => P(7)(281));
U_F8282: entity F port map(lamdaA => P(8)(282),lamdaB => P(8)(286),lamdaOut => P(7)(282));
U_F8283: entity F port map(lamdaA => P(8)(283),lamdaB => P(8)(287),lamdaOut => P(7)(283));
U_G8284: entity G port map(lamdaA => P(8)(280),lamdaB => P(8)(284),s => s(8)(140),lamdaOut => P(7)(284));
U_G8285: entity G port map(lamdaA => P(8)(281),lamdaB => P(8)(285),s => s(8)(141),lamdaOut => P(7)(285));
U_G8286: entity G port map(lamdaA => P(8)(282),lamdaB => P(8)(286),s => s(8)(142),lamdaOut => P(7)(286));
U_G8287: entity G port map(lamdaA => P(8)(283),lamdaB => P(8)(287),s => s(8)(143),lamdaOut => P(7)(287));
U_F8288: entity F port map(lamdaA => P(8)(288),lamdaB => P(8)(292),lamdaOut => P(7)(288));
U_F8289: entity F port map(lamdaA => P(8)(289),lamdaB => P(8)(293),lamdaOut => P(7)(289));
U_F8290: entity F port map(lamdaA => P(8)(290),lamdaB => P(8)(294),lamdaOut => P(7)(290));
U_F8291: entity F port map(lamdaA => P(8)(291),lamdaB => P(8)(295),lamdaOut => P(7)(291));
U_G8292: entity G port map(lamdaA => P(8)(288),lamdaB => P(8)(292),s => s(8)(144),lamdaOut => P(7)(292));
U_G8293: entity G port map(lamdaA => P(8)(289),lamdaB => P(8)(293),s => s(8)(145),lamdaOut => P(7)(293));
U_G8294: entity G port map(lamdaA => P(8)(290),lamdaB => P(8)(294),s => s(8)(146),lamdaOut => P(7)(294));
U_G8295: entity G port map(lamdaA => P(8)(291),lamdaB => P(8)(295),s => s(8)(147),lamdaOut => P(7)(295));
U_F8296: entity F port map(lamdaA => P(8)(296),lamdaB => P(8)(300),lamdaOut => P(7)(296));
U_F8297: entity F port map(lamdaA => P(8)(297),lamdaB => P(8)(301),lamdaOut => P(7)(297));
U_F8298: entity F port map(lamdaA => P(8)(298),lamdaB => P(8)(302),lamdaOut => P(7)(298));
U_F8299: entity F port map(lamdaA => P(8)(299),lamdaB => P(8)(303),lamdaOut => P(7)(299));
U_G8300: entity G port map(lamdaA => P(8)(296),lamdaB => P(8)(300),s => s(8)(148),lamdaOut => P(7)(300));
U_G8301: entity G port map(lamdaA => P(8)(297),lamdaB => P(8)(301),s => s(8)(149),lamdaOut => P(7)(301));
U_G8302: entity G port map(lamdaA => P(8)(298),lamdaB => P(8)(302),s => s(8)(150),lamdaOut => P(7)(302));
U_G8303: entity G port map(lamdaA => P(8)(299),lamdaB => P(8)(303),s => s(8)(151),lamdaOut => P(7)(303));
U_F8304: entity F port map(lamdaA => P(8)(304),lamdaB => P(8)(308),lamdaOut => P(7)(304));
U_F8305: entity F port map(lamdaA => P(8)(305),lamdaB => P(8)(309),lamdaOut => P(7)(305));
U_F8306: entity F port map(lamdaA => P(8)(306),lamdaB => P(8)(310),lamdaOut => P(7)(306));
U_F8307: entity F port map(lamdaA => P(8)(307),lamdaB => P(8)(311),lamdaOut => P(7)(307));
U_G8308: entity G port map(lamdaA => P(8)(304),lamdaB => P(8)(308),s => s(8)(152),lamdaOut => P(7)(308));
U_G8309: entity G port map(lamdaA => P(8)(305),lamdaB => P(8)(309),s => s(8)(153),lamdaOut => P(7)(309));
U_G8310: entity G port map(lamdaA => P(8)(306),lamdaB => P(8)(310),s => s(8)(154),lamdaOut => P(7)(310));
U_G8311: entity G port map(lamdaA => P(8)(307),lamdaB => P(8)(311),s => s(8)(155),lamdaOut => P(7)(311));
U_F8312: entity F port map(lamdaA => P(8)(312),lamdaB => P(8)(316),lamdaOut => P(7)(312));
U_F8313: entity F port map(lamdaA => P(8)(313),lamdaB => P(8)(317),lamdaOut => P(7)(313));
U_F8314: entity F port map(lamdaA => P(8)(314),lamdaB => P(8)(318),lamdaOut => P(7)(314));
U_F8315: entity F port map(lamdaA => P(8)(315),lamdaB => P(8)(319),lamdaOut => P(7)(315));
U_G8316: entity G port map(lamdaA => P(8)(312),lamdaB => P(8)(316),s => s(8)(156),lamdaOut => P(7)(316));
U_G8317: entity G port map(lamdaA => P(8)(313),lamdaB => P(8)(317),s => s(8)(157),lamdaOut => P(7)(317));
U_G8318: entity G port map(lamdaA => P(8)(314),lamdaB => P(8)(318),s => s(8)(158),lamdaOut => P(7)(318));
U_G8319: entity G port map(lamdaA => P(8)(315),lamdaB => P(8)(319),s => s(8)(159),lamdaOut => P(7)(319));
U_F8320: entity F port map(lamdaA => P(8)(320),lamdaB => P(8)(324),lamdaOut => P(7)(320));
U_F8321: entity F port map(lamdaA => P(8)(321),lamdaB => P(8)(325),lamdaOut => P(7)(321));
U_F8322: entity F port map(lamdaA => P(8)(322),lamdaB => P(8)(326),lamdaOut => P(7)(322));
U_F8323: entity F port map(lamdaA => P(8)(323),lamdaB => P(8)(327),lamdaOut => P(7)(323));
U_G8324: entity G port map(lamdaA => P(8)(320),lamdaB => P(8)(324),s => s(8)(160),lamdaOut => P(7)(324));
U_G8325: entity G port map(lamdaA => P(8)(321),lamdaB => P(8)(325),s => s(8)(161),lamdaOut => P(7)(325));
U_G8326: entity G port map(lamdaA => P(8)(322),lamdaB => P(8)(326),s => s(8)(162),lamdaOut => P(7)(326));
U_G8327: entity G port map(lamdaA => P(8)(323),lamdaB => P(8)(327),s => s(8)(163),lamdaOut => P(7)(327));
U_F8328: entity F port map(lamdaA => P(8)(328),lamdaB => P(8)(332),lamdaOut => P(7)(328));
U_F8329: entity F port map(lamdaA => P(8)(329),lamdaB => P(8)(333),lamdaOut => P(7)(329));
U_F8330: entity F port map(lamdaA => P(8)(330),lamdaB => P(8)(334),lamdaOut => P(7)(330));
U_F8331: entity F port map(lamdaA => P(8)(331),lamdaB => P(8)(335),lamdaOut => P(7)(331));
U_G8332: entity G port map(lamdaA => P(8)(328),lamdaB => P(8)(332),s => s(8)(164),lamdaOut => P(7)(332));
U_G8333: entity G port map(lamdaA => P(8)(329),lamdaB => P(8)(333),s => s(8)(165),lamdaOut => P(7)(333));
U_G8334: entity G port map(lamdaA => P(8)(330),lamdaB => P(8)(334),s => s(8)(166),lamdaOut => P(7)(334));
U_G8335: entity G port map(lamdaA => P(8)(331),lamdaB => P(8)(335),s => s(8)(167),lamdaOut => P(7)(335));
U_F8336: entity F port map(lamdaA => P(8)(336),lamdaB => P(8)(340),lamdaOut => P(7)(336));
U_F8337: entity F port map(lamdaA => P(8)(337),lamdaB => P(8)(341),lamdaOut => P(7)(337));
U_F8338: entity F port map(lamdaA => P(8)(338),lamdaB => P(8)(342),lamdaOut => P(7)(338));
U_F8339: entity F port map(lamdaA => P(8)(339),lamdaB => P(8)(343),lamdaOut => P(7)(339));
U_G8340: entity G port map(lamdaA => P(8)(336),lamdaB => P(8)(340),s => s(8)(168),lamdaOut => P(7)(340));
U_G8341: entity G port map(lamdaA => P(8)(337),lamdaB => P(8)(341),s => s(8)(169),lamdaOut => P(7)(341));
U_G8342: entity G port map(lamdaA => P(8)(338),lamdaB => P(8)(342),s => s(8)(170),lamdaOut => P(7)(342));
U_G8343: entity G port map(lamdaA => P(8)(339),lamdaB => P(8)(343),s => s(8)(171),lamdaOut => P(7)(343));
U_F8344: entity F port map(lamdaA => P(8)(344),lamdaB => P(8)(348),lamdaOut => P(7)(344));
U_F8345: entity F port map(lamdaA => P(8)(345),lamdaB => P(8)(349),lamdaOut => P(7)(345));
U_F8346: entity F port map(lamdaA => P(8)(346),lamdaB => P(8)(350),lamdaOut => P(7)(346));
U_F8347: entity F port map(lamdaA => P(8)(347),lamdaB => P(8)(351),lamdaOut => P(7)(347));
U_G8348: entity G port map(lamdaA => P(8)(344),lamdaB => P(8)(348),s => s(8)(172),lamdaOut => P(7)(348));
U_G8349: entity G port map(lamdaA => P(8)(345),lamdaB => P(8)(349),s => s(8)(173),lamdaOut => P(7)(349));
U_G8350: entity G port map(lamdaA => P(8)(346),lamdaB => P(8)(350),s => s(8)(174),lamdaOut => P(7)(350));
U_G8351: entity G port map(lamdaA => P(8)(347),lamdaB => P(8)(351),s => s(8)(175),lamdaOut => P(7)(351));
U_F8352: entity F port map(lamdaA => P(8)(352),lamdaB => P(8)(356),lamdaOut => P(7)(352));
U_F8353: entity F port map(lamdaA => P(8)(353),lamdaB => P(8)(357),lamdaOut => P(7)(353));
U_F8354: entity F port map(lamdaA => P(8)(354),lamdaB => P(8)(358),lamdaOut => P(7)(354));
U_F8355: entity F port map(lamdaA => P(8)(355),lamdaB => P(8)(359),lamdaOut => P(7)(355));
U_G8356: entity G port map(lamdaA => P(8)(352),lamdaB => P(8)(356),s => s(8)(176),lamdaOut => P(7)(356));
U_G8357: entity G port map(lamdaA => P(8)(353),lamdaB => P(8)(357),s => s(8)(177),lamdaOut => P(7)(357));
U_G8358: entity G port map(lamdaA => P(8)(354),lamdaB => P(8)(358),s => s(8)(178),lamdaOut => P(7)(358));
U_G8359: entity G port map(lamdaA => P(8)(355),lamdaB => P(8)(359),s => s(8)(179),lamdaOut => P(7)(359));
U_F8360: entity F port map(lamdaA => P(8)(360),lamdaB => P(8)(364),lamdaOut => P(7)(360));
U_F8361: entity F port map(lamdaA => P(8)(361),lamdaB => P(8)(365),lamdaOut => P(7)(361));
U_F8362: entity F port map(lamdaA => P(8)(362),lamdaB => P(8)(366),lamdaOut => P(7)(362));
U_F8363: entity F port map(lamdaA => P(8)(363),lamdaB => P(8)(367),lamdaOut => P(7)(363));
U_G8364: entity G port map(lamdaA => P(8)(360),lamdaB => P(8)(364),s => s(8)(180),lamdaOut => P(7)(364));
U_G8365: entity G port map(lamdaA => P(8)(361),lamdaB => P(8)(365),s => s(8)(181),lamdaOut => P(7)(365));
U_G8366: entity G port map(lamdaA => P(8)(362),lamdaB => P(8)(366),s => s(8)(182),lamdaOut => P(7)(366));
U_G8367: entity G port map(lamdaA => P(8)(363),lamdaB => P(8)(367),s => s(8)(183),lamdaOut => P(7)(367));
U_F8368: entity F port map(lamdaA => P(8)(368),lamdaB => P(8)(372),lamdaOut => P(7)(368));
U_F8369: entity F port map(lamdaA => P(8)(369),lamdaB => P(8)(373),lamdaOut => P(7)(369));
U_F8370: entity F port map(lamdaA => P(8)(370),lamdaB => P(8)(374),lamdaOut => P(7)(370));
U_F8371: entity F port map(lamdaA => P(8)(371),lamdaB => P(8)(375),lamdaOut => P(7)(371));
U_G8372: entity G port map(lamdaA => P(8)(368),lamdaB => P(8)(372),s => s(8)(184),lamdaOut => P(7)(372));
U_G8373: entity G port map(lamdaA => P(8)(369),lamdaB => P(8)(373),s => s(8)(185),lamdaOut => P(7)(373));
U_G8374: entity G port map(lamdaA => P(8)(370),lamdaB => P(8)(374),s => s(8)(186),lamdaOut => P(7)(374));
U_G8375: entity G port map(lamdaA => P(8)(371),lamdaB => P(8)(375),s => s(8)(187),lamdaOut => P(7)(375));
U_F8376: entity F port map(lamdaA => P(8)(376),lamdaB => P(8)(380),lamdaOut => P(7)(376));
U_F8377: entity F port map(lamdaA => P(8)(377),lamdaB => P(8)(381),lamdaOut => P(7)(377));
U_F8378: entity F port map(lamdaA => P(8)(378),lamdaB => P(8)(382),lamdaOut => P(7)(378));
U_F8379: entity F port map(lamdaA => P(8)(379),lamdaB => P(8)(383),lamdaOut => P(7)(379));
U_G8380: entity G port map(lamdaA => P(8)(376),lamdaB => P(8)(380),s => s(8)(188),lamdaOut => P(7)(380));
U_G8381: entity G port map(lamdaA => P(8)(377),lamdaB => P(8)(381),s => s(8)(189),lamdaOut => P(7)(381));
U_G8382: entity G port map(lamdaA => P(8)(378),lamdaB => P(8)(382),s => s(8)(190),lamdaOut => P(7)(382));
U_G8383: entity G port map(lamdaA => P(8)(379),lamdaB => P(8)(383),s => s(8)(191),lamdaOut => P(7)(383));
U_F8384: entity F port map(lamdaA => P(8)(384),lamdaB => P(8)(388),lamdaOut => P(7)(384));
U_F8385: entity F port map(lamdaA => P(8)(385),lamdaB => P(8)(389),lamdaOut => P(7)(385));
U_F8386: entity F port map(lamdaA => P(8)(386),lamdaB => P(8)(390),lamdaOut => P(7)(386));
U_F8387: entity F port map(lamdaA => P(8)(387),lamdaB => P(8)(391),lamdaOut => P(7)(387));
U_G8388: entity G port map(lamdaA => P(8)(384),lamdaB => P(8)(388),s => s(8)(192),lamdaOut => P(7)(388));
U_G8389: entity G port map(lamdaA => P(8)(385),lamdaB => P(8)(389),s => s(8)(193),lamdaOut => P(7)(389));
U_G8390: entity G port map(lamdaA => P(8)(386),lamdaB => P(8)(390),s => s(8)(194),lamdaOut => P(7)(390));
U_G8391: entity G port map(lamdaA => P(8)(387),lamdaB => P(8)(391),s => s(8)(195),lamdaOut => P(7)(391));
U_F8392: entity F port map(lamdaA => P(8)(392),lamdaB => P(8)(396),lamdaOut => P(7)(392));
U_F8393: entity F port map(lamdaA => P(8)(393),lamdaB => P(8)(397),lamdaOut => P(7)(393));
U_F8394: entity F port map(lamdaA => P(8)(394),lamdaB => P(8)(398),lamdaOut => P(7)(394));
U_F8395: entity F port map(lamdaA => P(8)(395),lamdaB => P(8)(399),lamdaOut => P(7)(395));
U_G8396: entity G port map(lamdaA => P(8)(392),lamdaB => P(8)(396),s => s(8)(196),lamdaOut => P(7)(396));
U_G8397: entity G port map(lamdaA => P(8)(393),lamdaB => P(8)(397),s => s(8)(197),lamdaOut => P(7)(397));
U_G8398: entity G port map(lamdaA => P(8)(394),lamdaB => P(8)(398),s => s(8)(198),lamdaOut => P(7)(398));
U_G8399: entity G port map(lamdaA => P(8)(395),lamdaB => P(8)(399),s => s(8)(199),lamdaOut => P(7)(399));
U_F8400: entity F port map(lamdaA => P(8)(400),lamdaB => P(8)(404),lamdaOut => P(7)(400));
U_F8401: entity F port map(lamdaA => P(8)(401),lamdaB => P(8)(405),lamdaOut => P(7)(401));
U_F8402: entity F port map(lamdaA => P(8)(402),lamdaB => P(8)(406),lamdaOut => P(7)(402));
U_F8403: entity F port map(lamdaA => P(8)(403),lamdaB => P(8)(407),lamdaOut => P(7)(403));
U_G8404: entity G port map(lamdaA => P(8)(400),lamdaB => P(8)(404),s => s(8)(200),lamdaOut => P(7)(404));
U_G8405: entity G port map(lamdaA => P(8)(401),lamdaB => P(8)(405),s => s(8)(201),lamdaOut => P(7)(405));
U_G8406: entity G port map(lamdaA => P(8)(402),lamdaB => P(8)(406),s => s(8)(202),lamdaOut => P(7)(406));
U_G8407: entity G port map(lamdaA => P(8)(403),lamdaB => P(8)(407),s => s(8)(203),lamdaOut => P(7)(407));
U_F8408: entity F port map(lamdaA => P(8)(408),lamdaB => P(8)(412),lamdaOut => P(7)(408));
U_F8409: entity F port map(lamdaA => P(8)(409),lamdaB => P(8)(413),lamdaOut => P(7)(409));
U_F8410: entity F port map(lamdaA => P(8)(410),lamdaB => P(8)(414),lamdaOut => P(7)(410));
U_F8411: entity F port map(lamdaA => P(8)(411),lamdaB => P(8)(415),lamdaOut => P(7)(411));
U_G8412: entity G port map(lamdaA => P(8)(408),lamdaB => P(8)(412),s => s(8)(204),lamdaOut => P(7)(412));
U_G8413: entity G port map(lamdaA => P(8)(409),lamdaB => P(8)(413),s => s(8)(205),lamdaOut => P(7)(413));
U_G8414: entity G port map(lamdaA => P(8)(410),lamdaB => P(8)(414),s => s(8)(206),lamdaOut => P(7)(414));
U_G8415: entity G port map(lamdaA => P(8)(411),lamdaB => P(8)(415),s => s(8)(207),lamdaOut => P(7)(415));
U_F8416: entity F port map(lamdaA => P(8)(416),lamdaB => P(8)(420),lamdaOut => P(7)(416));
U_F8417: entity F port map(lamdaA => P(8)(417),lamdaB => P(8)(421),lamdaOut => P(7)(417));
U_F8418: entity F port map(lamdaA => P(8)(418),lamdaB => P(8)(422),lamdaOut => P(7)(418));
U_F8419: entity F port map(lamdaA => P(8)(419),lamdaB => P(8)(423),lamdaOut => P(7)(419));
U_G8420: entity G port map(lamdaA => P(8)(416),lamdaB => P(8)(420),s => s(8)(208),lamdaOut => P(7)(420));
U_G8421: entity G port map(lamdaA => P(8)(417),lamdaB => P(8)(421),s => s(8)(209),lamdaOut => P(7)(421));
U_G8422: entity G port map(lamdaA => P(8)(418),lamdaB => P(8)(422),s => s(8)(210),lamdaOut => P(7)(422));
U_G8423: entity G port map(lamdaA => P(8)(419),lamdaB => P(8)(423),s => s(8)(211),lamdaOut => P(7)(423));
U_F8424: entity F port map(lamdaA => P(8)(424),lamdaB => P(8)(428),lamdaOut => P(7)(424));
U_F8425: entity F port map(lamdaA => P(8)(425),lamdaB => P(8)(429),lamdaOut => P(7)(425));
U_F8426: entity F port map(lamdaA => P(8)(426),lamdaB => P(8)(430),lamdaOut => P(7)(426));
U_F8427: entity F port map(lamdaA => P(8)(427),lamdaB => P(8)(431),lamdaOut => P(7)(427));
U_G8428: entity G port map(lamdaA => P(8)(424),lamdaB => P(8)(428),s => s(8)(212),lamdaOut => P(7)(428));
U_G8429: entity G port map(lamdaA => P(8)(425),lamdaB => P(8)(429),s => s(8)(213),lamdaOut => P(7)(429));
U_G8430: entity G port map(lamdaA => P(8)(426),lamdaB => P(8)(430),s => s(8)(214),lamdaOut => P(7)(430));
U_G8431: entity G port map(lamdaA => P(8)(427),lamdaB => P(8)(431),s => s(8)(215),lamdaOut => P(7)(431));
U_F8432: entity F port map(lamdaA => P(8)(432),lamdaB => P(8)(436),lamdaOut => P(7)(432));
U_F8433: entity F port map(lamdaA => P(8)(433),lamdaB => P(8)(437),lamdaOut => P(7)(433));
U_F8434: entity F port map(lamdaA => P(8)(434),lamdaB => P(8)(438),lamdaOut => P(7)(434));
U_F8435: entity F port map(lamdaA => P(8)(435),lamdaB => P(8)(439),lamdaOut => P(7)(435));
U_G8436: entity G port map(lamdaA => P(8)(432),lamdaB => P(8)(436),s => s(8)(216),lamdaOut => P(7)(436));
U_G8437: entity G port map(lamdaA => P(8)(433),lamdaB => P(8)(437),s => s(8)(217),lamdaOut => P(7)(437));
U_G8438: entity G port map(lamdaA => P(8)(434),lamdaB => P(8)(438),s => s(8)(218),lamdaOut => P(7)(438));
U_G8439: entity G port map(lamdaA => P(8)(435),lamdaB => P(8)(439),s => s(8)(219),lamdaOut => P(7)(439));
U_F8440: entity F port map(lamdaA => P(8)(440),lamdaB => P(8)(444),lamdaOut => P(7)(440));
U_F8441: entity F port map(lamdaA => P(8)(441),lamdaB => P(8)(445),lamdaOut => P(7)(441));
U_F8442: entity F port map(lamdaA => P(8)(442),lamdaB => P(8)(446),lamdaOut => P(7)(442));
U_F8443: entity F port map(lamdaA => P(8)(443),lamdaB => P(8)(447),lamdaOut => P(7)(443));
U_G8444: entity G port map(lamdaA => P(8)(440),lamdaB => P(8)(444),s => s(8)(220),lamdaOut => P(7)(444));
U_G8445: entity G port map(lamdaA => P(8)(441),lamdaB => P(8)(445),s => s(8)(221),lamdaOut => P(7)(445));
U_G8446: entity G port map(lamdaA => P(8)(442),lamdaB => P(8)(446),s => s(8)(222),lamdaOut => P(7)(446));
U_G8447: entity G port map(lamdaA => P(8)(443),lamdaB => P(8)(447),s => s(8)(223),lamdaOut => P(7)(447));
U_F8448: entity F port map(lamdaA => P(8)(448),lamdaB => P(8)(452),lamdaOut => P(7)(448));
U_F8449: entity F port map(lamdaA => P(8)(449),lamdaB => P(8)(453),lamdaOut => P(7)(449));
U_F8450: entity F port map(lamdaA => P(8)(450),lamdaB => P(8)(454),lamdaOut => P(7)(450));
U_F8451: entity F port map(lamdaA => P(8)(451),lamdaB => P(8)(455),lamdaOut => P(7)(451));
U_G8452: entity G port map(lamdaA => P(8)(448),lamdaB => P(8)(452),s => s(8)(224),lamdaOut => P(7)(452));
U_G8453: entity G port map(lamdaA => P(8)(449),lamdaB => P(8)(453),s => s(8)(225),lamdaOut => P(7)(453));
U_G8454: entity G port map(lamdaA => P(8)(450),lamdaB => P(8)(454),s => s(8)(226),lamdaOut => P(7)(454));
U_G8455: entity G port map(lamdaA => P(8)(451),lamdaB => P(8)(455),s => s(8)(227),lamdaOut => P(7)(455));
U_F8456: entity F port map(lamdaA => P(8)(456),lamdaB => P(8)(460),lamdaOut => P(7)(456));
U_F8457: entity F port map(lamdaA => P(8)(457),lamdaB => P(8)(461),lamdaOut => P(7)(457));
U_F8458: entity F port map(lamdaA => P(8)(458),lamdaB => P(8)(462),lamdaOut => P(7)(458));
U_F8459: entity F port map(lamdaA => P(8)(459),lamdaB => P(8)(463),lamdaOut => P(7)(459));
U_G8460: entity G port map(lamdaA => P(8)(456),lamdaB => P(8)(460),s => s(8)(228),lamdaOut => P(7)(460));
U_G8461: entity G port map(lamdaA => P(8)(457),lamdaB => P(8)(461),s => s(8)(229),lamdaOut => P(7)(461));
U_G8462: entity G port map(lamdaA => P(8)(458),lamdaB => P(8)(462),s => s(8)(230),lamdaOut => P(7)(462));
U_G8463: entity G port map(lamdaA => P(8)(459),lamdaB => P(8)(463),s => s(8)(231),lamdaOut => P(7)(463));
U_F8464: entity F port map(lamdaA => P(8)(464),lamdaB => P(8)(468),lamdaOut => P(7)(464));
U_F8465: entity F port map(lamdaA => P(8)(465),lamdaB => P(8)(469),lamdaOut => P(7)(465));
U_F8466: entity F port map(lamdaA => P(8)(466),lamdaB => P(8)(470),lamdaOut => P(7)(466));
U_F8467: entity F port map(lamdaA => P(8)(467),lamdaB => P(8)(471),lamdaOut => P(7)(467));
U_G8468: entity G port map(lamdaA => P(8)(464),lamdaB => P(8)(468),s => s(8)(232),lamdaOut => P(7)(468));
U_G8469: entity G port map(lamdaA => P(8)(465),lamdaB => P(8)(469),s => s(8)(233),lamdaOut => P(7)(469));
U_G8470: entity G port map(lamdaA => P(8)(466),lamdaB => P(8)(470),s => s(8)(234),lamdaOut => P(7)(470));
U_G8471: entity G port map(lamdaA => P(8)(467),lamdaB => P(8)(471),s => s(8)(235),lamdaOut => P(7)(471));
U_F8472: entity F port map(lamdaA => P(8)(472),lamdaB => P(8)(476),lamdaOut => P(7)(472));
U_F8473: entity F port map(lamdaA => P(8)(473),lamdaB => P(8)(477),lamdaOut => P(7)(473));
U_F8474: entity F port map(lamdaA => P(8)(474),lamdaB => P(8)(478),lamdaOut => P(7)(474));
U_F8475: entity F port map(lamdaA => P(8)(475),lamdaB => P(8)(479),lamdaOut => P(7)(475));
U_G8476: entity G port map(lamdaA => P(8)(472),lamdaB => P(8)(476),s => s(8)(236),lamdaOut => P(7)(476));
U_G8477: entity G port map(lamdaA => P(8)(473),lamdaB => P(8)(477),s => s(8)(237),lamdaOut => P(7)(477));
U_G8478: entity G port map(lamdaA => P(8)(474),lamdaB => P(8)(478),s => s(8)(238),lamdaOut => P(7)(478));
U_G8479: entity G port map(lamdaA => P(8)(475),lamdaB => P(8)(479),s => s(8)(239),lamdaOut => P(7)(479));
U_F8480: entity F port map(lamdaA => P(8)(480),lamdaB => P(8)(484),lamdaOut => P(7)(480));
U_F8481: entity F port map(lamdaA => P(8)(481),lamdaB => P(8)(485),lamdaOut => P(7)(481));
U_F8482: entity F port map(lamdaA => P(8)(482),lamdaB => P(8)(486),lamdaOut => P(7)(482));
U_F8483: entity F port map(lamdaA => P(8)(483),lamdaB => P(8)(487),lamdaOut => P(7)(483));
U_G8484: entity G port map(lamdaA => P(8)(480),lamdaB => P(8)(484),s => s(8)(240),lamdaOut => P(7)(484));
U_G8485: entity G port map(lamdaA => P(8)(481),lamdaB => P(8)(485),s => s(8)(241),lamdaOut => P(7)(485));
U_G8486: entity G port map(lamdaA => P(8)(482),lamdaB => P(8)(486),s => s(8)(242),lamdaOut => P(7)(486));
U_G8487: entity G port map(lamdaA => P(8)(483),lamdaB => P(8)(487),s => s(8)(243),lamdaOut => P(7)(487));
U_F8488: entity F port map(lamdaA => P(8)(488),lamdaB => P(8)(492),lamdaOut => P(7)(488));
U_F8489: entity F port map(lamdaA => P(8)(489),lamdaB => P(8)(493),lamdaOut => P(7)(489));
U_F8490: entity F port map(lamdaA => P(8)(490),lamdaB => P(8)(494),lamdaOut => P(7)(490));
U_F8491: entity F port map(lamdaA => P(8)(491),lamdaB => P(8)(495),lamdaOut => P(7)(491));
U_G8492: entity G port map(lamdaA => P(8)(488),lamdaB => P(8)(492),s => s(8)(244),lamdaOut => P(7)(492));
U_G8493: entity G port map(lamdaA => P(8)(489),lamdaB => P(8)(493),s => s(8)(245),lamdaOut => P(7)(493));
U_G8494: entity G port map(lamdaA => P(8)(490),lamdaB => P(8)(494),s => s(8)(246),lamdaOut => P(7)(494));
U_G8495: entity G port map(lamdaA => P(8)(491),lamdaB => P(8)(495),s => s(8)(247),lamdaOut => P(7)(495));
U_F8496: entity F port map(lamdaA => P(8)(496),lamdaB => P(8)(500),lamdaOut => P(7)(496));
U_F8497: entity F port map(lamdaA => P(8)(497),lamdaB => P(8)(501),lamdaOut => P(7)(497));
U_F8498: entity F port map(lamdaA => P(8)(498),lamdaB => P(8)(502),lamdaOut => P(7)(498));
U_F8499: entity F port map(lamdaA => P(8)(499),lamdaB => P(8)(503),lamdaOut => P(7)(499));
U_G8500: entity G port map(lamdaA => P(8)(496),lamdaB => P(8)(500),s => s(8)(248),lamdaOut => P(7)(500));
U_G8501: entity G port map(lamdaA => P(8)(497),lamdaB => P(8)(501),s => s(8)(249),lamdaOut => P(7)(501));
U_G8502: entity G port map(lamdaA => P(8)(498),lamdaB => P(8)(502),s => s(8)(250),lamdaOut => P(7)(502));
U_G8503: entity G port map(lamdaA => P(8)(499),lamdaB => P(8)(503),s => s(8)(251),lamdaOut => P(7)(503));
U_F8504: entity F port map(lamdaA => P(8)(504),lamdaB => P(8)(508),lamdaOut => P(7)(504));
U_F8505: entity F port map(lamdaA => P(8)(505),lamdaB => P(8)(509),lamdaOut => P(7)(505));
U_F8506: entity F port map(lamdaA => P(8)(506),lamdaB => P(8)(510),lamdaOut => P(7)(506));
U_F8507: entity F port map(lamdaA => P(8)(507),lamdaB => P(8)(511),lamdaOut => P(7)(507));
U_G8508: entity G port map(lamdaA => P(8)(504),lamdaB => P(8)(508),s => s(8)(252),lamdaOut => P(7)(508));
U_G8509: entity G port map(lamdaA => P(8)(505),lamdaB => P(8)(509),s => s(8)(253),lamdaOut => P(7)(509));
U_G8510: entity G port map(lamdaA => P(8)(506),lamdaB => P(8)(510),s => s(8)(254),lamdaOut => P(7)(510));
U_G8511: entity G port map(lamdaA => P(8)(507),lamdaB => P(8)(511),s => s(8)(255),lamdaOut => P(7)(511));
U_F8512: entity F port map(lamdaA => P(8)(512),lamdaB => P(8)(516),lamdaOut => P(7)(512));
U_F8513: entity F port map(lamdaA => P(8)(513),lamdaB => P(8)(517),lamdaOut => P(7)(513));
U_F8514: entity F port map(lamdaA => P(8)(514),lamdaB => P(8)(518),lamdaOut => P(7)(514));
U_F8515: entity F port map(lamdaA => P(8)(515),lamdaB => P(8)(519),lamdaOut => P(7)(515));
U_G8516: entity G port map(lamdaA => P(8)(512),lamdaB => P(8)(516),s => s(8)(256),lamdaOut => P(7)(516));
U_G8517: entity G port map(lamdaA => P(8)(513),lamdaB => P(8)(517),s => s(8)(257),lamdaOut => P(7)(517));
U_G8518: entity G port map(lamdaA => P(8)(514),lamdaB => P(8)(518),s => s(8)(258),lamdaOut => P(7)(518));
U_G8519: entity G port map(lamdaA => P(8)(515),lamdaB => P(8)(519),s => s(8)(259),lamdaOut => P(7)(519));
U_F8520: entity F port map(lamdaA => P(8)(520),lamdaB => P(8)(524),lamdaOut => P(7)(520));
U_F8521: entity F port map(lamdaA => P(8)(521),lamdaB => P(8)(525),lamdaOut => P(7)(521));
U_F8522: entity F port map(lamdaA => P(8)(522),lamdaB => P(8)(526),lamdaOut => P(7)(522));
U_F8523: entity F port map(lamdaA => P(8)(523),lamdaB => P(8)(527),lamdaOut => P(7)(523));
U_G8524: entity G port map(lamdaA => P(8)(520),lamdaB => P(8)(524),s => s(8)(260),lamdaOut => P(7)(524));
U_G8525: entity G port map(lamdaA => P(8)(521),lamdaB => P(8)(525),s => s(8)(261),lamdaOut => P(7)(525));
U_G8526: entity G port map(lamdaA => P(8)(522),lamdaB => P(8)(526),s => s(8)(262),lamdaOut => P(7)(526));
U_G8527: entity G port map(lamdaA => P(8)(523),lamdaB => P(8)(527),s => s(8)(263),lamdaOut => P(7)(527));
U_F8528: entity F port map(lamdaA => P(8)(528),lamdaB => P(8)(532),lamdaOut => P(7)(528));
U_F8529: entity F port map(lamdaA => P(8)(529),lamdaB => P(8)(533),lamdaOut => P(7)(529));
U_F8530: entity F port map(lamdaA => P(8)(530),lamdaB => P(8)(534),lamdaOut => P(7)(530));
U_F8531: entity F port map(lamdaA => P(8)(531),lamdaB => P(8)(535),lamdaOut => P(7)(531));
U_G8532: entity G port map(lamdaA => P(8)(528),lamdaB => P(8)(532),s => s(8)(264),lamdaOut => P(7)(532));
U_G8533: entity G port map(lamdaA => P(8)(529),lamdaB => P(8)(533),s => s(8)(265),lamdaOut => P(7)(533));
U_G8534: entity G port map(lamdaA => P(8)(530),lamdaB => P(8)(534),s => s(8)(266),lamdaOut => P(7)(534));
U_G8535: entity G port map(lamdaA => P(8)(531),lamdaB => P(8)(535),s => s(8)(267),lamdaOut => P(7)(535));
U_F8536: entity F port map(lamdaA => P(8)(536),lamdaB => P(8)(540),lamdaOut => P(7)(536));
U_F8537: entity F port map(lamdaA => P(8)(537),lamdaB => P(8)(541),lamdaOut => P(7)(537));
U_F8538: entity F port map(lamdaA => P(8)(538),lamdaB => P(8)(542),lamdaOut => P(7)(538));
U_F8539: entity F port map(lamdaA => P(8)(539),lamdaB => P(8)(543),lamdaOut => P(7)(539));
U_G8540: entity G port map(lamdaA => P(8)(536),lamdaB => P(8)(540),s => s(8)(268),lamdaOut => P(7)(540));
U_G8541: entity G port map(lamdaA => P(8)(537),lamdaB => P(8)(541),s => s(8)(269),lamdaOut => P(7)(541));
U_G8542: entity G port map(lamdaA => P(8)(538),lamdaB => P(8)(542),s => s(8)(270),lamdaOut => P(7)(542));
U_G8543: entity G port map(lamdaA => P(8)(539),lamdaB => P(8)(543),s => s(8)(271),lamdaOut => P(7)(543));
U_F8544: entity F port map(lamdaA => P(8)(544),lamdaB => P(8)(548),lamdaOut => P(7)(544));
U_F8545: entity F port map(lamdaA => P(8)(545),lamdaB => P(8)(549),lamdaOut => P(7)(545));
U_F8546: entity F port map(lamdaA => P(8)(546),lamdaB => P(8)(550),lamdaOut => P(7)(546));
U_F8547: entity F port map(lamdaA => P(8)(547),lamdaB => P(8)(551),lamdaOut => P(7)(547));
U_G8548: entity G port map(lamdaA => P(8)(544),lamdaB => P(8)(548),s => s(8)(272),lamdaOut => P(7)(548));
U_G8549: entity G port map(lamdaA => P(8)(545),lamdaB => P(8)(549),s => s(8)(273),lamdaOut => P(7)(549));
U_G8550: entity G port map(lamdaA => P(8)(546),lamdaB => P(8)(550),s => s(8)(274),lamdaOut => P(7)(550));
U_G8551: entity G port map(lamdaA => P(8)(547),lamdaB => P(8)(551),s => s(8)(275),lamdaOut => P(7)(551));
U_F8552: entity F port map(lamdaA => P(8)(552),lamdaB => P(8)(556),lamdaOut => P(7)(552));
U_F8553: entity F port map(lamdaA => P(8)(553),lamdaB => P(8)(557),lamdaOut => P(7)(553));
U_F8554: entity F port map(lamdaA => P(8)(554),lamdaB => P(8)(558),lamdaOut => P(7)(554));
U_F8555: entity F port map(lamdaA => P(8)(555),lamdaB => P(8)(559),lamdaOut => P(7)(555));
U_G8556: entity G port map(lamdaA => P(8)(552),lamdaB => P(8)(556),s => s(8)(276),lamdaOut => P(7)(556));
U_G8557: entity G port map(lamdaA => P(8)(553),lamdaB => P(8)(557),s => s(8)(277),lamdaOut => P(7)(557));
U_G8558: entity G port map(lamdaA => P(8)(554),lamdaB => P(8)(558),s => s(8)(278),lamdaOut => P(7)(558));
U_G8559: entity G port map(lamdaA => P(8)(555),lamdaB => P(8)(559),s => s(8)(279),lamdaOut => P(7)(559));
U_F8560: entity F port map(lamdaA => P(8)(560),lamdaB => P(8)(564),lamdaOut => P(7)(560));
U_F8561: entity F port map(lamdaA => P(8)(561),lamdaB => P(8)(565),lamdaOut => P(7)(561));
U_F8562: entity F port map(lamdaA => P(8)(562),lamdaB => P(8)(566),lamdaOut => P(7)(562));
U_F8563: entity F port map(lamdaA => P(8)(563),lamdaB => P(8)(567),lamdaOut => P(7)(563));
U_G8564: entity G port map(lamdaA => P(8)(560),lamdaB => P(8)(564),s => s(8)(280),lamdaOut => P(7)(564));
U_G8565: entity G port map(lamdaA => P(8)(561),lamdaB => P(8)(565),s => s(8)(281),lamdaOut => P(7)(565));
U_G8566: entity G port map(lamdaA => P(8)(562),lamdaB => P(8)(566),s => s(8)(282),lamdaOut => P(7)(566));
U_G8567: entity G port map(lamdaA => P(8)(563),lamdaB => P(8)(567),s => s(8)(283),lamdaOut => P(7)(567));
U_F8568: entity F port map(lamdaA => P(8)(568),lamdaB => P(8)(572),lamdaOut => P(7)(568));
U_F8569: entity F port map(lamdaA => P(8)(569),lamdaB => P(8)(573),lamdaOut => P(7)(569));
U_F8570: entity F port map(lamdaA => P(8)(570),lamdaB => P(8)(574),lamdaOut => P(7)(570));
U_F8571: entity F port map(lamdaA => P(8)(571),lamdaB => P(8)(575),lamdaOut => P(7)(571));
U_G8572: entity G port map(lamdaA => P(8)(568),lamdaB => P(8)(572),s => s(8)(284),lamdaOut => P(7)(572));
U_G8573: entity G port map(lamdaA => P(8)(569),lamdaB => P(8)(573),s => s(8)(285),lamdaOut => P(7)(573));
U_G8574: entity G port map(lamdaA => P(8)(570),lamdaB => P(8)(574),s => s(8)(286),lamdaOut => P(7)(574));
U_G8575: entity G port map(lamdaA => P(8)(571),lamdaB => P(8)(575),s => s(8)(287),lamdaOut => P(7)(575));
U_F8576: entity F port map(lamdaA => P(8)(576),lamdaB => P(8)(580),lamdaOut => P(7)(576));
U_F8577: entity F port map(lamdaA => P(8)(577),lamdaB => P(8)(581),lamdaOut => P(7)(577));
U_F8578: entity F port map(lamdaA => P(8)(578),lamdaB => P(8)(582),lamdaOut => P(7)(578));
U_F8579: entity F port map(lamdaA => P(8)(579),lamdaB => P(8)(583),lamdaOut => P(7)(579));
U_G8580: entity G port map(lamdaA => P(8)(576),lamdaB => P(8)(580),s => s(8)(288),lamdaOut => P(7)(580));
U_G8581: entity G port map(lamdaA => P(8)(577),lamdaB => P(8)(581),s => s(8)(289),lamdaOut => P(7)(581));
U_G8582: entity G port map(lamdaA => P(8)(578),lamdaB => P(8)(582),s => s(8)(290),lamdaOut => P(7)(582));
U_G8583: entity G port map(lamdaA => P(8)(579),lamdaB => P(8)(583),s => s(8)(291),lamdaOut => P(7)(583));
U_F8584: entity F port map(lamdaA => P(8)(584),lamdaB => P(8)(588),lamdaOut => P(7)(584));
U_F8585: entity F port map(lamdaA => P(8)(585),lamdaB => P(8)(589),lamdaOut => P(7)(585));
U_F8586: entity F port map(lamdaA => P(8)(586),lamdaB => P(8)(590),lamdaOut => P(7)(586));
U_F8587: entity F port map(lamdaA => P(8)(587),lamdaB => P(8)(591),lamdaOut => P(7)(587));
U_G8588: entity G port map(lamdaA => P(8)(584),lamdaB => P(8)(588),s => s(8)(292),lamdaOut => P(7)(588));
U_G8589: entity G port map(lamdaA => P(8)(585),lamdaB => P(8)(589),s => s(8)(293),lamdaOut => P(7)(589));
U_G8590: entity G port map(lamdaA => P(8)(586),lamdaB => P(8)(590),s => s(8)(294),lamdaOut => P(7)(590));
U_G8591: entity G port map(lamdaA => P(8)(587),lamdaB => P(8)(591),s => s(8)(295),lamdaOut => P(7)(591));
U_F8592: entity F port map(lamdaA => P(8)(592),lamdaB => P(8)(596),lamdaOut => P(7)(592));
U_F8593: entity F port map(lamdaA => P(8)(593),lamdaB => P(8)(597),lamdaOut => P(7)(593));
U_F8594: entity F port map(lamdaA => P(8)(594),lamdaB => P(8)(598),lamdaOut => P(7)(594));
U_F8595: entity F port map(lamdaA => P(8)(595),lamdaB => P(8)(599),lamdaOut => P(7)(595));
U_G8596: entity G port map(lamdaA => P(8)(592),lamdaB => P(8)(596),s => s(8)(296),lamdaOut => P(7)(596));
U_G8597: entity G port map(lamdaA => P(8)(593),lamdaB => P(8)(597),s => s(8)(297),lamdaOut => P(7)(597));
U_G8598: entity G port map(lamdaA => P(8)(594),lamdaB => P(8)(598),s => s(8)(298),lamdaOut => P(7)(598));
U_G8599: entity G port map(lamdaA => P(8)(595),lamdaB => P(8)(599),s => s(8)(299),lamdaOut => P(7)(599));
U_F8600: entity F port map(lamdaA => P(8)(600),lamdaB => P(8)(604),lamdaOut => P(7)(600));
U_F8601: entity F port map(lamdaA => P(8)(601),lamdaB => P(8)(605),lamdaOut => P(7)(601));
U_F8602: entity F port map(lamdaA => P(8)(602),lamdaB => P(8)(606),lamdaOut => P(7)(602));
U_F8603: entity F port map(lamdaA => P(8)(603),lamdaB => P(8)(607),lamdaOut => P(7)(603));
U_G8604: entity G port map(lamdaA => P(8)(600),lamdaB => P(8)(604),s => s(8)(300),lamdaOut => P(7)(604));
U_G8605: entity G port map(lamdaA => P(8)(601),lamdaB => P(8)(605),s => s(8)(301),lamdaOut => P(7)(605));
U_G8606: entity G port map(lamdaA => P(8)(602),lamdaB => P(8)(606),s => s(8)(302),lamdaOut => P(7)(606));
U_G8607: entity G port map(lamdaA => P(8)(603),lamdaB => P(8)(607),s => s(8)(303),lamdaOut => P(7)(607));
U_F8608: entity F port map(lamdaA => P(8)(608),lamdaB => P(8)(612),lamdaOut => P(7)(608));
U_F8609: entity F port map(lamdaA => P(8)(609),lamdaB => P(8)(613),lamdaOut => P(7)(609));
U_F8610: entity F port map(lamdaA => P(8)(610),lamdaB => P(8)(614),lamdaOut => P(7)(610));
U_F8611: entity F port map(lamdaA => P(8)(611),lamdaB => P(8)(615),lamdaOut => P(7)(611));
U_G8612: entity G port map(lamdaA => P(8)(608),lamdaB => P(8)(612),s => s(8)(304),lamdaOut => P(7)(612));
U_G8613: entity G port map(lamdaA => P(8)(609),lamdaB => P(8)(613),s => s(8)(305),lamdaOut => P(7)(613));
U_G8614: entity G port map(lamdaA => P(8)(610),lamdaB => P(8)(614),s => s(8)(306),lamdaOut => P(7)(614));
U_G8615: entity G port map(lamdaA => P(8)(611),lamdaB => P(8)(615),s => s(8)(307),lamdaOut => P(7)(615));
U_F8616: entity F port map(lamdaA => P(8)(616),lamdaB => P(8)(620),lamdaOut => P(7)(616));
U_F8617: entity F port map(lamdaA => P(8)(617),lamdaB => P(8)(621),lamdaOut => P(7)(617));
U_F8618: entity F port map(lamdaA => P(8)(618),lamdaB => P(8)(622),lamdaOut => P(7)(618));
U_F8619: entity F port map(lamdaA => P(8)(619),lamdaB => P(8)(623),lamdaOut => P(7)(619));
U_G8620: entity G port map(lamdaA => P(8)(616),lamdaB => P(8)(620),s => s(8)(308),lamdaOut => P(7)(620));
U_G8621: entity G port map(lamdaA => P(8)(617),lamdaB => P(8)(621),s => s(8)(309),lamdaOut => P(7)(621));
U_G8622: entity G port map(lamdaA => P(8)(618),lamdaB => P(8)(622),s => s(8)(310),lamdaOut => P(7)(622));
U_G8623: entity G port map(lamdaA => P(8)(619),lamdaB => P(8)(623),s => s(8)(311),lamdaOut => P(7)(623));
U_F8624: entity F port map(lamdaA => P(8)(624),lamdaB => P(8)(628),lamdaOut => P(7)(624));
U_F8625: entity F port map(lamdaA => P(8)(625),lamdaB => P(8)(629),lamdaOut => P(7)(625));
U_F8626: entity F port map(lamdaA => P(8)(626),lamdaB => P(8)(630),lamdaOut => P(7)(626));
U_F8627: entity F port map(lamdaA => P(8)(627),lamdaB => P(8)(631),lamdaOut => P(7)(627));
U_G8628: entity G port map(lamdaA => P(8)(624),lamdaB => P(8)(628),s => s(8)(312),lamdaOut => P(7)(628));
U_G8629: entity G port map(lamdaA => P(8)(625),lamdaB => P(8)(629),s => s(8)(313),lamdaOut => P(7)(629));
U_G8630: entity G port map(lamdaA => P(8)(626),lamdaB => P(8)(630),s => s(8)(314),lamdaOut => P(7)(630));
U_G8631: entity G port map(lamdaA => P(8)(627),lamdaB => P(8)(631),s => s(8)(315),lamdaOut => P(7)(631));
U_F8632: entity F port map(lamdaA => P(8)(632),lamdaB => P(8)(636),lamdaOut => P(7)(632));
U_F8633: entity F port map(lamdaA => P(8)(633),lamdaB => P(8)(637),lamdaOut => P(7)(633));
U_F8634: entity F port map(lamdaA => P(8)(634),lamdaB => P(8)(638),lamdaOut => P(7)(634));
U_F8635: entity F port map(lamdaA => P(8)(635),lamdaB => P(8)(639),lamdaOut => P(7)(635));
U_G8636: entity G port map(lamdaA => P(8)(632),lamdaB => P(8)(636),s => s(8)(316),lamdaOut => P(7)(636));
U_G8637: entity G port map(lamdaA => P(8)(633),lamdaB => P(8)(637),s => s(8)(317),lamdaOut => P(7)(637));
U_G8638: entity G port map(lamdaA => P(8)(634),lamdaB => P(8)(638),s => s(8)(318),lamdaOut => P(7)(638));
U_G8639: entity G port map(lamdaA => P(8)(635),lamdaB => P(8)(639),s => s(8)(319),lamdaOut => P(7)(639));
U_F8640: entity F port map(lamdaA => P(8)(640),lamdaB => P(8)(644),lamdaOut => P(7)(640));
U_F8641: entity F port map(lamdaA => P(8)(641),lamdaB => P(8)(645),lamdaOut => P(7)(641));
U_F8642: entity F port map(lamdaA => P(8)(642),lamdaB => P(8)(646),lamdaOut => P(7)(642));
U_F8643: entity F port map(lamdaA => P(8)(643),lamdaB => P(8)(647),lamdaOut => P(7)(643));
U_G8644: entity G port map(lamdaA => P(8)(640),lamdaB => P(8)(644),s => s(8)(320),lamdaOut => P(7)(644));
U_G8645: entity G port map(lamdaA => P(8)(641),lamdaB => P(8)(645),s => s(8)(321),lamdaOut => P(7)(645));
U_G8646: entity G port map(lamdaA => P(8)(642),lamdaB => P(8)(646),s => s(8)(322),lamdaOut => P(7)(646));
U_G8647: entity G port map(lamdaA => P(8)(643),lamdaB => P(8)(647),s => s(8)(323),lamdaOut => P(7)(647));
U_F8648: entity F port map(lamdaA => P(8)(648),lamdaB => P(8)(652),lamdaOut => P(7)(648));
U_F8649: entity F port map(lamdaA => P(8)(649),lamdaB => P(8)(653),lamdaOut => P(7)(649));
U_F8650: entity F port map(lamdaA => P(8)(650),lamdaB => P(8)(654),lamdaOut => P(7)(650));
U_F8651: entity F port map(lamdaA => P(8)(651),lamdaB => P(8)(655),lamdaOut => P(7)(651));
U_G8652: entity G port map(lamdaA => P(8)(648),lamdaB => P(8)(652),s => s(8)(324),lamdaOut => P(7)(652));
U_G8653: entity G port map(lamdaA => P(8)(649),lamdaB => P(8)(653),s => s(8)(325),lamdaOut => P(7)(653));
U_G8654: entity G port map(lamdaA => P(8)(650),lamdaB => P(8)(654),s => s(8)(326),lamdaOut => P(7)(654));
U_G8655: entity G port map(lamdaA => P(8)(651),lamdaB => P(8)(655),s => s(8)(327),lamdaOut => P(7)(655));
U_F8656: entity F port map(lamdaA => P(8)(656),lamdaB => P(8)(660),lamdaOut => P(7)(656));
U_F8657: entity F port map(lamdaA => P(8)(657),lamdaB => P(8)(661),lamdaOut => P(7)(657));
U_F8658: entity F port map(lamdaA => P(8)(658),lamdaB => P(8)(662),lamdaOut => P(7)(658));
U_F8659: entity F port map(lamdaA => P(8)(659),lamdaB => P(8)(663),lamdaOut => P(7)(659));
U_G8660: entity G port map(lamdaA => P(8)(656),lamdaB => P(8)(660),s => s(8)(328),lamdaOut => P(7)(660));
U_G8661: entity G port map(lamdaA => P(8)(657),lamdaB => P(8)(661),s => s(8)(329),lamdaOut => P(7)(661));
U_G8662: entity G port map(lamdaA => P(8)(658),lamdaB => P(8)(662),s => s(8)(330),lamdaOut => P(7)(662));
U_G8663: entity G port map(lamdaA => P(8)(659),lamdaB => P(8)(663),s => s(8)(331),lamdaOut => P(7)(663));
U_F8664: entity F port map(lamdaA => P(8)(664),lamdaB => P(8)(668),lamdaOut => P(7)(664));
U_F8665: entity F port map(lamdaA => P(8)(665),lamdaB => P(8)(669),lamdaOut => P(7)(665));
U_F8666: entity F port map(lamdaA => P(8)(666),lamdaB => P(8)(670),lamdaOut => P(7)(666));
U_F8667: entity F port map(lamdaA => P(8)(667),lamdaB => P(8)(671),lamdaOut => P(7)(667));
U_G8668: entity G port map(lamdaA => P(8)(664),lamdaB => P(8)(668),s => s(8)(332),lamdaOut => P(7)(668));
U_G8669: entity G port map(lamdaA => P(8)(665),lamdaB => P(8)(669),s => s(8)(333),lamdaOut => P(7)(669));
U_G8670: entity G port map(lamdaA => P(8)(666),lamdaB => P(8)(670),s => s(8)(334),lamdaOut => P(7)(670));
U_G8671: entity G port map(lamdaA => P(8)(667),lamdaB => P(8)(671),s => s(8)(335),lamdaOut => P(7)(671));
U_F8672: entity F port map(lamdaA => P(8)(672),lamdaB => P(8)(676),lamdaOut => P(7)(672));
U_F8673: entity F port map(lamdaA => P(8)(673),lamdaB => P(8)(677),lamdaOut => P(7)(673));
U_F8674: entity F port map(lamdaA => P(8)(674),lamdaB => P(8)(678),lamdaOut => P(7)(674));
U_F8675: entity F port map(lamdaA => P(8)(675),lamdaB => P(8)(679),lamdaOut => P(7)(675));
U_G8676: entity G port map(lamdaA => P(8)(672),lamdaB => P(8)(676),s => s(8)(336),lamdaOut => P(7)(676));
U_G8677: entity G port map(lamdaA => P(8)(673),lamdaB => P(8)(677),s => s(8)(337),lamdaOut => P(7)(677));
U_G8678: entity G port map(lamdaA => P(8)(674),lamdaB => P(8)(678),s => s(8)(338),lamdaOut => P(7)(678));
U_G8679: entity G port map(lamdaA => P(8)(675),lamdaB => P(8)(679),s => s(8)(339),lamdaOut => P(7)(679));
U_F8680: entity F port map(lamdaA => P(8)(680),lamdaB => P(8)(684),lamdaOut => P(7)(680));
U_F8681: entity F port map(lamdaA => P(8)(681),lamdaB => P(8)(685),lamdaOut => P(7)(681));
U_F8682: entity F port map(lamdaA => P(8)(682),lamdaB => P(8)(686),lamdaOut => P(7)(682));
U_F8683: entity F port map(lamdaA => P(8)(683),lamdaB => P(8)(687),lamdaOut => P(7)(683));
U_G8684: entity G port map(lamdaA => P(8)(680),lamdaB => P(8)(684),s => s(8)(340),lamdaOut => P(7)(684));
U_G8685: entity G port map(lamdaA => P(8)(681),lamdaB => P(8)(685),s => s(8)(341),lamdaOut => P(7)(685));
U_G8686: entity G port map(lamdaA => P(8)(682),lamdaB => P(8)(686),s => s(8)(342),lamdaOut => P(7)(686));
U_G8687: entity G port map(lamdaA => P(8)(683),lamdaB => P(8)(687),s => s(8)(343),lamdaOut => P(7)(687));
U_F8688: entity F port map(lamdaA => P(8)(688),lamdaB => P(8)(692),lamdaOut => P(7)(688));
U_F8689: entity F port map(lamdaA => P(8)(689),lamdaB => P(8)(693),lamdaOut => P(7)(689));
U_F8690: entity F port map(lamdaA => P(8)(690),lamdaB => P(8)(694),lamdaOut => P(7)(690));
U_F8691: entity F port map(lamdaA => P(8)(691),lamdaB => P(8)(695),lamdaOut => P(7)(691));
U_G8692: entity G port map(lamdaA => P(8)(688),lamdaB => P(8)(692),s => s(8)(344),lamdaOut => P(7)(692));
U_G8693: entity G port map(lamdaA => P(8)(689),lamdaB => P(8)(693),s => s(8)(345),lamdaOut => P(7)(693));
U_G8694: entity G port map(lamdaA => P(8)(690),lamdaB => P(8)(694),s => s(8)(346),lamdaOut => P(7)(694));
U_G8695: entity G port map(lamdaA => P(8)(691),lamdaB => P(8)(695),s => s(8)(347),lamdaOut => P(7)(695));
U_F8696: entity F port map(lamdaA => P(8)(696),lamdaB => P(8)(700),lamdaOut => P(7)(696));
U_F8697: entity F port map(lamdaA => P(8)(697),lamdaB => P(8)(701),lamdaOut => P(7)(697));
U_F8698: entity F port map(lamdaA => P(8)(698),lamdaB => P(8)(702),lamdaOut => P(7)(698));
U_F8699: entity F port map(lamdaA => P(8)(699),lamdaB => P(8)(703),lamdaOut => P(7)(699));
U_G8700: entity G port map(lamdaA => P(8)(696),lamdaB => P(8)(700),s => s(8)(348),lamdaOut => P(7)(700));
U_G8701: entity G port map(lamdaA => P(8)(697),lamdaB => P(8)(701),s => s(8)(349),lamdaOut => P(7)(701));
U_G8702: entity G port map(lamdaA => P(8)(698),lamdaB => P(8)(702),s => s(8)(350),lamdaOut => P(7)(702));
U_G8703: entity G port map(lamdaA => P(8)(699),lamdaB => P(8)(703),s => s(8)(351),lamdaOut => P(7)(703));
U_F8704: entity F port map(lamdaA => P(8)(704),lamdaB => P(8)(708),lamdaOut => P(7)(704));
U_F8705: entity F port map(lamdaA => P(8)(705),lamdaB => P(8)(709),lamdaOut => P(7)(705));
U_F8706: entity F port map(lamdaA => P(8)(706),lamdaB => P(8)(710),lamdaOut => P(7)(706));
U_F8707: entity F port map(lamdaA => P(8)(707),lamdaB => P(8)(711),lamdaOut => P(7)(707));
U_G8708: entity G port map(lamdaA => P(8)(704),lamdaB => P(8)(708),s => s(8)(352),lamdaOut => P(7)(708));
U_G8709: entity G port map(lamdaA => P(8)(705),lamdaB => P(8)(709),s => s(8)(353),lamdaOut => P(7)(709));
U_G8710: entity G port map(lamdaA => P(8)(706),lamdaB => P(8)(710),s => s(8)(354),lamdaOut => P(7)(710));
U_G8711: entity G port map(lamdaA => P(8)(707),lamdaB => P(8)(711),s => s(8)(355),lamdaOut => P(7)(711));
U_F8712: entity F port map(lamdaA => P(8)(712),lamdaB => P(8)(716),lamdaOut => P(7)(712));
U_F8713: entity F port map(lamdaA => P(8)(713),lamdaB => P(8)(717),lamdaOut => P(7)(713));
U_F8714: entity F port map(lamdaA => P(8)(714),lamdaB => P(8)(718),lamdaOut => P(7)(714));
U_F8715: entity F port map(lamdaA => P(8)(715),lamdaB => P(8)(719),lamdaOut => P(7)(715));
U_G8716: entity G port map(lamdaA => P(8)(712),lamdaB => P(8)(716),s => s(8)(356),lamdaOut => P(7)(716));
U_G8717: entity G port map(lamdaA => P(8)(713),lamdaB => P(8)(717),s => s(8)(357),lamdaOut => P(7)(717));
U_G8718: entity G port map(lamdaA => P(8)(714),lamdaB => P(8)(718),s => s(8)(358),lamdaOut => P(7)(718));
U_G8719: entity G port map(lamdaA => P(8)(715),lamdaB => P(8)(719),s => s(8)(359),lamdaOut => P(7)(719));
U_F8720: entity F port map(lamdaA => P(8)(720),lamdaB => P(8)(724),lamdaOut => P(7)(720));
U_F8721: entity F port map(lamdaA => P(8)(721),lamdaB => P(8)(725),lamdaOut => P(7)(721));
U_F8722: entity F port map(lamdaA => P(8)(722),lamdaB => P(8)(726),lamdaOut => P(7)(722));
U_F8723: entity F port map(lamdaA => P(8)(723),lamdaB => P(8)(727),lamdaOut => P(7)(723));
U_G8724: entity G port map(lamdaA => P(8)(720),lamdaB => P(8)(724),s => s(8)(360),lamdaOut => P(7)(724));
U_G8725: entity G port map(lamdaA => P(8)(721),lamdaB => P(8)(725),s => s(8)(361),lamdaOut => P(7)(725));
U_G8726: entity G port map(lamdaA => P(8)(722),lamdaB => P(8)(726),s => s(8)(362),lamdaOut => P(7)(726));
U_G8727: entity G port map(lamdaA => P(8)(723),lamdaB => P(8)(727),s => s(8)(363),lamdaOut => P(7)(727));
U_F8728: entity F port map(lamdaA => P(8)(728),lamdaB => P(8)(732),lamdaOut => P(7)(728));
U_F8729: entity F port map(lamdaA => P(8)(729),lamdaB => P(8)(733),lamdaOut => P(7)(729));
U_F8730: entity F port map(lamdaA => P(8)(730),lamdaB => P(8)(734),lamdaOut => P(7)(730));
U_F8731: entity F port map(lamdaA => P(8)(731),lamdaB => P(8)(735),lamdaOut => P(7)(731));
U_G8732: entity G port map(lamdaA => P(8)(728),lamdaB => P(8)(732),s => s(8)(364),lamdaOut => P(7)(732));
U_G8733: entity G port map(lamdaA => P(8)(729),lamdaB => P(8)(733),s => s(8)(365),lamdaOut => P(7)(733));
U_G8734: entity G port map(lamdaA => P(8)(730),lamdaB => P(8)(734),s => s(8)(366),lamdaOut => P(7)(734));
U_G8735: entity G port map(lamdaA => P(8)(731),lamdaB => P(8)(735),s => s(8)(367),lamdaOut => P(7)(735));
U_F8736: entity F port map(lamdaA => P(8)(736),lamdaB => P(8)(740),lamdaOut => P(7)(736));
U_F8737: entity F port map(lamdaA => P(8)(737),lamdaB => P(8)(741),lamdaOut => P(7)(737));
U_F8738: entity F port map(lamdaA => P(8)(738),lamdaB => P(8)(742),lamdaOut => P(7)(738));
U_F8739: entity F port map(lamdaA => P(8)(739),lamdaB => P(8)(743),lamdaOut => P(7)(739));
U_G8740: entity G port map(lamdaA => P(8)(736),lamdaB => P(8)(740),s => s(8)(368),lamdaOut => P(7)(740));
U_G8741: entity G port map(lamdaA => P(8)(737),lamdaB => P(8)(741),s => s(8)(369),lamdaOut => P(7)(741));
U_G8742: entity G port map(lamdaA => P(8)(738),lamdaB => P(8)(742),s => s(8)(370),lamdaOut => P(7)(742));
U_G8743: entity G port map(lamdaA => P(8)(739),lamdaB => P(8)(743),s => s(8)(371),lamdaOut => P(7)(743));
U_F8744: entity F port map(lamdaA => P(8)(744),lamdaB => P(8)(748),lamdaOut => P(7)(744));
U_F8745: entity F port map(lamdaA => P(8)(745),lamdaB => P(8)(749),lamdaOut => P(7)(745));
U_F8746: entity F port map(lamdaA => P(8)(746),lamdaB => P(8)(750),lamdaOut => P(7)(746));
U_F8747: entity F port map(lamdaA => P(8)(747),lamdaB => P(8)(751),lamdaOut => P(7)(747));
U_G8748: entity G port map(lamdaA => P(8)(744),lamdaB => P(8)(748),s => s(8)(372),lamdaOut => P(7)(748));
U_G8749: entity G port map(lamdaA => P(8)(745),lamdaB => P(8)(749),s => s(8)(373),lamdaOut => P(7)(749));
U_G8750: entity G port map(lamdaA => P(8)(746),lamdaB => P(8)(750),s => s(8)(374),lamdaOut => P(7)(750));
U_G8751: entity G port map(lamdaA => P(8)(747),lamdaB => P(8)(751),s => s(8)(375),lamdaOut => P(7)(751));
U_F8752: entity F port map(lamdaA => P(8)(752),lamdaB => P(8)(756),lamdaOut => P(7)(752));
U_F8753: entity F port map(lamdaA => P(8)(753),lamdaB => P(8)(757),lamdaOut => P(7)(753));
U_F8754: entity F port map(lamdaA => P(8)(754),lamdaB => P(8)(758),lamdaOut => P(7)(754));
U_F8755: entity F port map(lamdaA => P(8)(755),lamdaB => P(8)(759),lamdaOut => P(7)(755));
U_G8756: entity G port map(lamdaA => P(8)(752),lamdaB => P(8)(756),s => s(8)(376),lamdaOut => P(7)(756));
U_G8757: entity G port map(lamdaA => P(8)(753),lamdaB => P(8)(757),s => s(8)(377),lamdaOut => P(7)(757));
U_G8758: entity G port map(lamdaA => P(8)(754),lamdaB => P(8)(758),s => s(8)(378),lamdaOut => P(7)(758));
U_G8759: entity G port map(lamdaA => P(8)(755),lamdaB => P(8)(759),s => s(8)(379),lamdaOut => P(7)(759));
U_F8760: entity F port map(lamdaA => P(8)(760),lamdaB => P(8)(764),lamdaOut => P(7)(760));
U_F8761: entity F port map(lamdaA => P(8)(761),lamdaB => P(8)(765),lamdaOut => P(7)(761));
U_F8762: entity F port map(lamdaA => P(8)(762),lamdaB => P(8)(766),lamdaOut => P(7)(762));
U_F8763: entity F port map(lamdaA => P(8)(763),lamdaB => P(8)(767),lamdaOut => P(7)(763));
U_G8764: entity G port map(lamdaA => P(8)(760),lamdaB => P(8)(764),s => s(8)(380),lamdaOut => P(7)(764));
U_G8765: entity G port map(lamdaA => P(8)(761),lamdaB => P(8)(765),s => s(8)(381),lamdaOut => P(7)(765));
U_G8766: entity G port map(lamdaA => P(8)(762),lamdaB => P(8)(766),s => s(8)(382),lamdaOut => P(7)(766));
U_G8767: entity G port map(lamdaA => P(8)(763),lamdaB => P(8)(767),s => s(8)(383),lamdaOut => P(7)(767));
U_F8768: entity F port map(lamdaA => P(8)(768),lamdaB => P(8)(772),lamdaOut => P(7)(768));
U_F8769: entity F port map(lamdaA => P(8)(769),lamdaB => P(8)(773),lamdaOut => P(7)(769));
U_F8770: entity F port map(lamdaA => P(8)(770),lamdaB => P(8)(774),lamdaOut => P(7)(770));
U_F8771: entity F port map(lamdaA => P(8)(771),lamdaB => P(8)(775),lamdaOut => P(7)(771));
U_G8772: entity G port map(lamdaA => P(8)(768),lamdaB => P(8)(772),s => s(8)(384),lamdaOut => P(7)(772));
U_G8773: entity G port map(lamdaA => P(8)(769),lamdaB => P(8)(773),s => s(8)(385),lamdaOut => P(7)(773));
U_G8774: entity G port map(lamdaA => P(8)(770),lamdaB => P(8)(774),s => s(8)(386),lamdaOut => P(7)(774));
U_G8775: entity G port map(lamdaA => P(8)(771),lamdaB => P(8)(775),s => s(8)(387),lamdaOut => P(7)(775));
U_F8776: entity F port map(lamdaA => P(8)(776),lamdaB => P(8)(780),lamdaOut => P(7)(776));
U_F8777: entity F port map(lamdaA => P(8)(777),lamdaB => P(8)(781),lamdaOut => P(7)(777));
U_F8778: entity F port map(lamdaA => P(8)(778),lamdaB => P(8)(782),lamdaOut => P(7)(778));
U_F8779: entity F port map(lamdaA => P(8)(779),lamdaB => P(8)(783),lamdaOut => P(7)(779));
U_G8780: entity G port map(lamdaA => P(8)(776),lamdaB => P(8)(780),s => s(8)(388),lamdaOut => P(7)(780));
U_G8781: entity G port map(lamdaA => P(8)(777),lamdaB => P(8)(781),s => s(8)(389),lamdaOut => P(7)(781));
U_G8782: entity G port map(lamdaA => P(8)(778),lamdaB => P(8)(782),s => s(8)(390),lamdaOut => P(7)(782));
U_G8783: entity G port map(lamdaA => P(8)(779),lamdaB => P(8)(783),s => s(8)(391),lamdaOut => P(7)(783));
U_F8784: entity F port map(lamdaA => P(8)(784),lamdaB => P(8)(788),lamdaOut => P(7)(784));
U_F8785: entity F port map(lamdaA => P(8)(785),lamdaB => P(8)(789),lamdaOut => P(7)(785));
U_F8786: entity F port map(lamdaA => P(8)(786),lamdaB => P(8)(790),lamdaOut => P(7)(786));
U_F8787: entity F port map(lamdaA => P(8)(787),lamdaB => P(8)(791),lamdaOut => P(7)(787));
U_G8788: entity G port map(lamdaA => P(8)(784),lamdaB => P(8)(788),s => s(8)(392),lamdaOut => P(7)(788));
U_G8789: entity G port map(lamdaA => P(8)(785),lamdaB => P(8)(789),s => s(8)(393),lamdaOut => P(7)(789));
U_G8790: entity G port map(lamdaA => P(8)(786),lamdaB => P(8)(790),s => s(8)(394),lamdaOut => P(7)(790));
U_G8791: entity G port map(lamdaA => P(8)(787),lamdaB => P(8)(791),s => s(8)(395),lamdaOut => P(7)(791));
U_F8792: entity F port map(lamdaA => P(8)(792),lamdaB => P(8)(796),lamdaOut => P(7)(792));
U_F8793: entity F port map(lamdaA => P(8)(793),lamdaB => P(8)(797),lamdaOut => P(7)(793));
U_F8794: entity F port map(lamdaA => P(8)(794),lamdaB => P(8)(798),lamdaOut => P(7)(794));
U_F8795: entity F port map(lamdaA => P(8)(795),lamdaB => P(8)(799),lamdaOut => P(7)(795));
U_G8796: entity G port map(lamdaA => P(8)(792),lamdaB => P(8)(796),s => s(8)(396),lamdaOut => P(7)(796));
U_G8797: entity G port map(lamdaA => P(8)(793),lamdaB => P(8)(797),s => s(8)(397),lamdaOut => P(7)(797));
U_G8798: entity G port map(lamdaA => P(8)(794),lamdaB => P(8)(798),s => s(8)(398),lamdaOut => P(7)(798));
U_G8799: entity G port map(lamdaA => P(8)(795),lamdaB => P(8)(799),s => s(8)(399),lamdaOut => P(7)(799));
U_F8800: entity F port map(lamdaA => P(8)(800),lamdaB => P(8)(804),lamdaOut => P(7)(800));
U_F8801: entity F port map(lamdaA => P(8)(801),lamdaB => P(8)(805),lamdaOut => P(7)(801));
U_F8802: entity F port map(lamdaA => P(8)(802),lamdaB => P(8)(806),lamdaOut => P(7)(802));
U_F8803: entity F port map(lamdaA => P(8)(803),lamdaB => P(8)(807),lamdaOut => P(7)(803));
U_G8804: entity G port map(lamdaA => P(8)(800),lamdaB => P(8)(804),s => s(8)(400),lamdaOut => P(7)(804));
U_G8805: entity G port map(lamdaA => P(8)(801),lamdaB => P(8)(805),s => s(8)(401),lamdaOut => P(7)(805));
U_G8806: entity G port map(lamdaA => P(8)(802),lamdaB => P(8)(806),s => s(8)(402),lamdaOut => P(7)(806));
U_G8807: entity G port map(lamdaA => P(8)(803),lamdaB => P(8)(807),s => s(8)(403),lamdaOut => P(7)(807));
U_F8808: entity F port map(lamdaA => P(8)(808),lamdaB => P(8)(812),lamdaOut => P(7)(808));
U_F8809: entity F port map(lamdaA => P(8)(809),lamdaB => P(8)(813),lamdaOut => P(7)(809));
U_F8810: entity F port map(lamdaA => P(8)(810),lamdaB => P(8)(814),lamdaOut => P(7)(810));
U_F8811: entity F port map(lamdaA => P(8)(811),lamdaB => P(8)(815),lamdaOut => P(7)(811));
U_G8812: entity G port map(lamdaA => P(8)(808),lamdaB => P(8)(812),s => s(8)(404),lamdaOut => P(7)(812));
U_G8813: entity G port map(lamdaA => P(8)(809),lamdaB => P(8)(813),s => s(8)(405),lamdaOut => P(7)(813));
U_G8814: entity G port map(lamdaA => P(8)(810),lamdaB => P(8)(814),s => s(8)(406),lamdaOut => P(7)(814));
U_G8815: entity G port map(lamdaA => P(8)(811),lamdaB => P(8)(815),s => s(8)(407),lamdaOut => P(7)(815));
U_F8816: entity F port map(lamdaA => P(8)(816),lamdaB => P(8)(820),lamdaOut => P(7)(816));
U_F8817: entity F port map(lamdaA => P(8)(817),lamdaB => P(8)(821),lamdaOut => P(7)(817));
U_F8818: entity F port map(lamdaA => P(8)(818),lamdaB => P(8)(822),lamdaOut => P(7)(818));
U_F8819: entity F port map(lamdaA => P(8)(819),lamdaB => P(8)(823),lamdaOut => P(7)(819));
U_G8820: entity G port map(lamdaA => P(8)(816),lamdaB => P(8)(820),s => s(8)(408),lamdaOut => P(7)(820));
U_G8821: entity G port map(lamdaA => P(8)(817),lamdaB => P(8)(821),s => s(8)(409),lamdaOut => P(7)(821));
U_G8822: entity G port map(lamdaA => P(8)(818),lamdaB => P(8)(822),s => s(8)(410),lamdaOut => P(7)(822));
U_G8823: entity G port map(lamdaA => P(8)(819),lamdaB => P(8)(823),s => s(8)(411),lamdaOut => P(7)(823));
U_F8824: entity F port map(lamdaA => P(8)(824),lamdaB => P(8)(828),lamdaOut => P(7)(824));
U_F8825: entity F port map(lamdaA => P(8)(825),lamdaB => P(8)(829),lamdaOut => P(7)(825));
U_F8826: entity F port map(lamdaA => P(8)(826),lamdaB => P(8)(830),lamdaOut => P(7)(826));
U_F8827: entity F port map(lamdaA => P(8)(827),lamdaB => P(8)(831),lamdaOut => P(7)(827));
U_G8828: entity G port map(lamdaA => P(8)(824),lamdaB => P(8)(828),s => s(8)(412),lamdaOut => P(7)(828));
U_G8829: entity G port map(lamdaA => P(8)(825),lamdaB => P(8)(829),s => s(8)(413),lamdaOut => P(7)(829));
U_G8830: entity G port map(lamdaA => P(8)(826),lamdaB => P(8)(830),s => s(8)(414),lamdaOut => P(7)(830));
U_G8831: entity G port map(lamdaA => P(8)(827),lamdaB => P(8)(831),s => s(8)(415),lamdaOut => P(7)(831));
U_F8832: entity F port map(lamdaA => P(8)(832),lamdaB => P(8)(836),lamdaOut => P(7)(832));
U_F8833: entity F port map(lamdaA => P(8)(833),lamdaB => P(8)(837),lamdaOut => P(7)(833));
U_F8834: entity F port map(lamdaA => P(8)(834),lamdaB => P(8)(838),lamdaOut => P(7)(834));
U_F8835: entity F port map(lamdaA => P(8)(835),lamdaB => P(8)(839),lamdaOut => P(7)(835));
U_G8836: entity G port map(lamdaA => P(8)(832),lamdaB => P(8)(836),s => s(8)(416),lamdaOut => P(7)(836));
U_G8837: entity G port map(lamdaA => P(8)(833),lamdaB => P(8)(837),s => s(8)(417),lamdaOut => P(7)(837));
U_G8838: entity G port map(lamdaA => P(8)(834),lamdaB => P(8)(838),s => s(8)(418),lamdaOut => P(7)(838));
U_G8839: entity G port map(lamdaA => P(8)(835),lamdaB => P(8)(839),s => s(8)(419),lamdaOut => P(7)(839));
U_F8840: entity F port map(lamdaA => P(8)(840),lamdaB => P(8)(844),lamdaOut => P(7)(840));
U_F8841: entity F port map(lamdaA => P(8)(841),lamdaB => P(8)(845),lamdaOut => P(7)(841));
U_F8842: entity F port map(lamdaA => P(8)(842),lamdaB => P(8)(846),lamdaOut => P(7)(842));
U_F8843: entity F port map(lamdaA => P(8)(843),lamdaB => P(8)(847),lamdaOut => P(7)(843));
U_G8844: entity G port map(lamdaA => P(8)(840),lamdaB => P(8)(844),s => s(8)(420),lamdaOut => P(7)(844));
U_G8845: entity G port map(lamdaA => P(8)(841),lamdaB => P(8)(845),s => s(8)(421),lamdaOut => P(7)(845));
U_G8846: entity G port map(lamdaA => P(8)(842),lamdaB => P(8)(846),s => s(8)(422),lamdaOut => P(7)(846));
U_G8847: entity G port map(lamdaA => P(8)(843),lamdaB => P(8)(847),s => s(8)(423),lamdaOut => P(7)(847));
U_F8848: entity F port map(lamdaA => P(8)(848),lamdaB => P(8)(852),lamdaOut => P(7)(848));
U_F8849: entity F port map(lamdaA => P(8)(849),lamdaB => P(8)(853),lamdaOut => P(7)(849));
U_F8850: entity F port map(lamdaA => P(8)(850),lamdaB => P(8)(854),lamdaOut => P(7)(850));
U_F8851: entity F port map(lamdaA => P(8)(851),lamdaB => P(8)(855),lamdaOut => P(7)(851));
U_G8852: entity G port map(lamdaA => P(8)(848),lamdaB => P(8)(852),s => s(8)(424),lamdaOut => P(7)(852));
U_G8853: entity G port map(lamdaA => P(8)(849),lamdaB => P(8)(853),s => s(8)(425),lamdaOut => P(7)(853));
U_G8854: entity G port map(lamdaA => P(8)(850),lamdaB => P(8)(854),s => s(8)(426),lamdaOut => P(7)(854));
U_G8855: entity G port map(lamdaA => P(8)(851),lamdaB => P(8)(855),s => s(8)(427),lamdaOut => P(7)(855));
U_F8856: entity F port map(lamdaA => P(8)(856),lamdaB => P(8)(860),lamdaOut => P(7)(856));
U_F8857: entity F port map(lamdaA => P(8)(857),lamdaB => P(8)(861),lamdaOut => P(7)(857));
U_F8858: entity F port map(lamdaA => P(8)(858),lamdaB => P(8)(862),lamdaOut => P(7)(858));
U_F8859: entity F port map(lamdaA => P(8)(859),lamdaB => P(8)(863),lamdaOut => P(7)(859));
U_G8860: entity G port map(lamdaA => P(8)(856),lamdaB => P(8)(860),s => s(8)(428),lamdaOut => P(7)(860));
U_G8861: entity G port map(lamdaA => P(8)(857),lamdaB => P(8)(861),s => s(8)(429),lamdaOut => P(7)(861));
U_G8862: entity G port map(lamdaA => P(8)(858),lamdaB => P(8)(862),s => s(8)(430),lamdaOut => P(7)(862));
U_G8863: entity G port map(lamdaA => P(8)(859),lamdaB => P(8)(863),s => s(8)(431),lamdaOut => P(7)(863));
U_F8864: entity F port map(lamdaA => P(8)(864),lamdaB => P(8)(868),lamdaOut => P(7)(864));
U_F8865: entity F port map(lamdaA => P(8)(865),lamdaB => P(8)(869),lamdaOut => P(7)(865));
U_F8866: entity F port map(lamdaA => P(8)(866),lamdaB => P(8)(870),lamdaOut => P(7)(866));
U_F8867: entity F port map(lamdaA => P(8)(867),lamdaB => P(8)(871),lamdaOut => P(7)(867));
U_G8868: entity G port map(lamdaA => P(8)(864),lamdaB => P(8)(868),s => s(8)(432),lamdaOut => P(7)(868));
U_G8869: entity G port map(lamdaA => P(8)(865),lamdaB => P(8)(869),s => s(8)(433),lamdaOut => P(7)(869));
U_G8870: entity G port map(lamdaA => P(8)(866),lamdaB => P(8)(870),s => s(8)(434),lamdaOut => P(7)(870));
U_G8871: entity G port map(lamdaA => P(8)(867),lamdaB => P(8)(871),s => s(8)(435),lamdaOut => P(7)(871));
U_F8872: entity F port map(lamdaA => P(8)(872),lamdaB => P(8)(876),lamdaOut => P(7)(872));
U_F8873: entity F port map(lamdaA => P(8)(873),lamdaB => P(8)(877),lamdaOut => P(7)(873));
U_F8874: entity F port map(lamdaA => P(8)(874),lamdaB => P(8)(878),lamdaOut => P(7)(874));
U_F8875: entity F port map(lamdaA => P(8)(875),lamdaB => P(8)(879),lamdaOut => P(7)(875));
U_G8876: entity G port map(lamdaA => P(8)(872),lamdaB => P(8)(876),s => s(8)(436),lamdaOut => P(7)(876));
U_G8877: entity G port map(lamdaA => P(8)(873),lamdaB => P(8)(877),s => s(8)(437),lamdaOut => P(7)(877));
U_G8878: entity G port map(lamdaA => P(8)(874),lamdaB => P(8)(878),s => s(8)(438),lamdaOut => P(7)(878));
U_G8879: entity G port map(lamdaA => P(8)(875),lamdaB => P(8)(879),s => s(8)(439),lamdaOut => P(7)(879));
U_F8880: entity F port map(lamdaA => P(8)(880),lamdaB => P(8)(884),lamdaOut => P(7)(880));
U_F8881: entity F port map(lamdaA => P(8)(881),lamdaB => P(8)(885),lamdaOut => P(7)(881));
U_F8882: entity F port map(lamdaA => P(8)(882),lamdaB => P(8)(886),lamdaOut => P(7)(882));
U_F8883: entity F port map(lamdaA => P(8)(883),lamdaB => P(8)(887),lamdaOut => P(7)(883));
U_G8884: entity G port map(lamdaA => P(8)(880),lamdaB => P(8)(884),s => s(8)(440),lamdaOut => P(7)(884));
U_G8885: entity G port map(lamdaA => P(8)(881),lamdaB => P(8)(885),s => s(8)(441),lamdaOut => P(7)(885));
U_G8886: entity G port map(lamdaA => P(8)(882),lamdaB => P(8)(886),s => s(8)(442),lamdaOut => P(7)(886));
U_G8887: entity G port map(lamdaA => P(8)(883),lamdaB => P(8)(887),s => s(8)(443),lamdaOut => P(7)(887));
U_F8888: entity F port map(lamdaA => P(8)(888),lamdaB => P(8)(892),lamdaOut => P(7)(888));
U_F8889: entity F port map(lamdaA => P(8)(889),lamdaB => P(8)(893),lamdaOut => P(7)(889));
U_F8890: entity F port map(lamdaA => P(8)(890),lamdaB => P(8)(894),lamdaOut => P(7)(890));
U_F8891: entity F port map(lamdaA => P(8)(891),lamdaB => P(8)(895),lamdaOut => P(7)(891));
U_G8892: entity G port map(lamdaA => P(8)(888),lamdaB => P(8)(892),s => s(8)(444),lamdaOut => P(7)(892));
U_G8893: entity G port map(lamdaA => P(8)(889),lamdaB => P(8)(893),s => s(8)(445),lamdaOut => P(7)(893));
U_G8894: entity G port map(lamdaA => P(8)(890),lamdaB => P(8)(894),s => s(8)(446),lamdaOut => P(7)(894));
U_G8895: entity G port map(lamdaA => P(8)(891),lamdaB => P(8)(895),s => s(8)(447),lamdaOut => P(7)(895));
U_F8896: entity F port map(lamdaA => P(8)(896),lamdaB => P(8)(900),lamdaOut => P(7)(896));
U_F8897: entity F port map(lamdaA => P(8)(897),lamdaB => P(8)(901),lamdaOut => P(7)(897));
U_F8898: entity F port map(lamdaA => P(8)(898),lamdaB => P(8)(902),lamdaOut => P(7)(898));
U_F8899: entity F port map(lamdaA => P(8)(899),lamdaB => P(8)(903),lamdaOut => P(7)(899));
U_G8900: entity G port map(lamdaA => P(8)(896),lamdaB => P(8)(900),s => s(8)(448),lamdaOut => P(7)(900));
U_G8901: entity G port map(lamdaA => P(8)(897),lamdaB => P(8)(901),s => s(8)(449),lamdaOut => P(7)(901));
U_G8902: entity G port map(lamdaA => P(8)(898),lamdaB => P(8)(902),s => s(8)(450),lamdaOut => P(7)(902));
U_G8903: entity G port map(lamdaA => P(8)(899),lamdaB => P(8)(903),s => s(8)(451),lamdaOut => P(7)(903));
U_F8904: entity F port map(lamdaA => P(8)(904),lamdaB => P(8)(908),lamdaOut => P(7)(904));
U_F8905: entity F port map(lamdaA => P(8)(905),lamdaB => P(8)(909),lamdaOut => P(7)(905));
U_F8906: entity F port map(lamdaA => P(8)(906),lamdaB => P(8)(910),lamdaOut => P(7)(906));
U_F8907: entity F port map(lamdaA => P(8)(907),lamdaB => P(8)(911),lamdaOut => P(7)(907));
U_G8908: entity G port map(lamdaA => P(8)(904),lamdaB => P(8)(908),s => s(8)(452),lamdaOut => P(7)(908));
U_G8909: entity G port map(lamdaA => P(8)(905),lamdaB => P(8)(909),s => s(8)(453),lamdaOut => P(7)(909));
U_G8910: entity G port map(lamdaA => P(8)(906),lamdaB => P(8)(910),s => s(8)(454),lamdaOut => P(7)(910));
U_G8911: entity G port map(lamdaA => P(8)(907),lamdaB => P(8)(911),s => s(8)(455),lamdaOut => P(7)(911));
U_F8912: entity F port map(lamdaA => P(8)(912),lamdaB => P(8)(916),lamdaOut => P(7)(912));
U_F8913: entity F port map(lamdaA => P(8)(913),lamdaB => P(8)(917),lamdaOut => P(7)(913));
U_F8914: entity F port map(lamdaA => P(8)(914),lamdaB => P(8)(918),lamdaOut => P(7)(914));
U_F8915: entity F port map(lamdaA => P(8)(915),lamdaB => P(8)(919),lamdaOut => P(7)(915));
U_G8916: entity G port map(lamdaA => P(8)(912),lamdaB => P(8)(916),s => s(8)(456),lamdaOut => P(7)(916));
U_G8917: entity G port map(lamdaA => P(8)(913),lamdaB => P(8)(917),s => s(8)(457),lamdaOut => P(7)(917));
U_G8918: entity G port map(lamdaA => P(8)(914),lamdaB => P(8)(918),s => s(8)(458),lamdaOut => P(7)(918));
U_G8919: entity G port map(lamdaA => P(8)(915),lamdaB => P(8)(919),s => s(8)(459),lamdaOut => P(7)(919));
U_F8920: entity F port map(lamdaA => P(8)(920),lamdaB => P(8)(924),lamdaOut => P(7)(920));
U_F8921: entity F port map(lamdaA => P(8)(921),lamdaB => P(8)(925),lamdaOut => P(7)(921));
U_F8922: entity F port map(lamdaA => P(8)(922),lamdaB => P(8)(926),lamdaOut => P(7)(922));
U_F8923: entity F port map(lamdaA => P(8)(923),lamdaB => P(8)(927),lamdaOut => P(7)(923));
U_G8924: entity G port map(lamdaA => P(8)(920),lamdaB => P(8)(924),s => s(8)(460),lamdaOut => P(7)(924));
U_G8925: entity G port map(lamdaA => P(8)(921),lamdaB => P(8)(925),s => s(8)(461),lamdaOut => P(7)(925));
U_G8926: entity G port map(lamdaA => P(8)(922),lamdaB => P(8)(926),s => s(8)(462),lamdaOut => P(7)(926));
U_G8927: entity G port map(lamdaA => P(8)(923),lamdaB => P(8)(927),s => s(8)(463),lamdaOut => P(7)(927));
U_F8928: entity F port map(lamdaA => P(8)(928),lamdaB => P(8)(932),lamdaOut => P(7)(928));
U_F8929: entity F port map(lamdaA => P(8)(929),lamdaB => P(8)(933),lamdaOut => P(7)(929));
U_F8930: entity F port map(lamdaA => P(8)(930),lamdaB => P(8)(934),lamdaOut => P(7)(930));
U_F8931: entity F port map(lamdaA => P(8)(931),lamdaB => P(8)(935),lamdaOut => P(7)(931));
U_G8932: entity G port map(lamdaA => P(8)(928),lamdaB => P(8)(932),s => s(8)(464),lamdaOut => P(7)(932));
U_G8933: entity G port map(lamdaA => P(8)(929),lamdaB => P(8)(933),s => s(8)(465),lamdaOut => P(7)(933));
U_G8934: entity G port map(lamdaA => P(8)(930),lamdaB => P(8)(934),s => s(8)(466),lamdaOut => P(7)(934));
U_G8935: entity G port map(lamdaA => P(8)(931),lamdaB => P(8)(935),s => s(8)(467),lamdaOut => P(7)(935));
U_F8936: entity F port map(lamdaA => P(8)(936),lamdaB => P(8)(940),lamdaOut => P(7)(936));
U_F8937: entity F port map(lamdaA => P(8)(937),lamdaB => P(8)(941),lamdaOut => P(7)(937));
U_F8938: entity F port map(lamdaA => P(8)(938),lamdaB => P(8)(942),lamdaOut => P(7)(938));
U_F8939: entity F port map(lamdaA => P(8)(939),lamdaB => P(8)(943),lamdaOut => P(7)(939));
U_G8940: entity G port map(lamdaA => P(8)(936),lamdaB => P(8)(940),s => s(8)(468),lamdaOut => P(7)(940));
U_G8941: entity G port map(lamdaA => P(8)(937),lamdaB => P(8)(941),s => s(8)(469),lamdaOut => P(7)(941));
U_G8942: entity G port map(lamdaA => P(8)(938),lamdaB => P(8)(942),s => s(8)(470),lamdaOut => P(7)(942));
U_G8943: entity G port map(lamdaA => P(8)(939),lamdaB => P(8)(943),s => s(8)(471),lamdaOut => P(7)(943));
U_F8944: entity F port map(lamdaA => P(8)(944),lamdaB => P(8)(948),lamdaOut => P(7)(944));
U_F8945: entity F port map(lamdaA => P(8)(945),lamdaB => P(8)(949),lamdaOut => P(7)(945));
U_F8946: entity F port map(lamdaA => P(8)(946),lamdaB => P(8)(950),lamdaOut => P(7)(946));
U_F8947: entity F port map(lamdaA => P(8)(947),lamdaB => P(8)(951),lamdaOut => P(7)(947));
U_G8948: entity G port map(lamdaA => P(8)(944),lamdaB => P(8)(948),s => s(8)(472),lamdaOut => P(7)(948));
U_G8949: entity G port map(lamdaA => P(8)(945),lamdaB => P(8)(949),s => s(8)(473),lamdaOut => P(7)(949));
U_G8950: entity G port map(lamdaA => P(8)(946),lamdaB => P(8)(950),s => s(8)(474),lamdaOut => P(7)(950));
U_G8951: entity G port map(lamdaA => P(8)(947),lamdaB => P(8)(951),s => s(8)(475),lamdaOut => P(7)(951));
U_F8952: entity F port map(lamdaA => P(8)(952),lamdaB => P(8)(956),lamdaOut => P(7)(952));
U_F8953: entity F port map(lamdaA => P(8)(953),lamdaB => P(8)(957),lamdaOut => P(7)(953));
U_F8954: entity F port map(lamdaA => P(8)(954),lamdaB => P(8)(958),lamdaOut => P(7)(954));
U_F8955: entity F port map(lamdaA => P(8)(955),lamdaB => P(8)(959),lamdaOut => P(7)(955));
U_G8956: entity G port map(lamdaA => P(8)(952),lamdaB => P(8)(956),s => s(8)(476),lamdaOut => P(7)(956));
U_G8957: entity G port map(lamdaA => P(8)(953),lamdaB => P(8)(957),s => s(8)(477),lamdaOut => P(7)(957));
U_G8958: entity G port map(lamdaA => P(8)(954),lamdaB => P(8)(958),s => s(8)(478),lamdaOut => P(7)(958));
U_G8959: entity G port map(lamdaA => P(8)(955),lamdaB => P(8)(959),s => s(8)(479),lamdaOut => P(7)(959));
U_F8960: entity F port map(lamdaA => P(8)(960),lamdaB => P(8)(964),lamdaOut => P(7)(960));
U_F8961: entity F port map(lamdaA => P(8)(961),lamdaB => P(8)(965),lamdaOut => P(7)(961));
U_F8962: entity F port map(lamdaA => P(8)(962),lamdaB => P(8)(966),lamdaOut => P(7)(962));
U_F8963: entity F port map(lamdaA => P(8)(963),lamdaB => P(8)(967),lamdaOut => P(7)(963));
U_G8964: entity G port map(lamdaA => P(8)(960),lamdaB => P(8)(964),s => s(8)(480),lamdaOut => P(7)(964));
U_G8965: entity G port map(lamdaA => P(8)(961),lamdaB => P(8)(965),s => s(8)(481),lamdaOut => P(7)(965));
U_G8966: entity G port map(lamdaA => P(8)(962),lamdaB => P(8)(966),s => s(8)(482),lamdaOut => P(7)(966));
U_G8967: entity G port map(lamdaA => P(8)(963),lamdaB => P(8)(967),s => s(8)(483),lamdaOut => P(7)(967));
U_F8968: entity F port map(lamdaA => P(8)(968),lamdaB => P(8)(972),lamdaOut => P(7)(968));
U_F8969: entity F port map(lamdaA => P(8)(969),lamdaB => P(8)(973),lamdaOut => P(7)(969));
U_F8970: entity F port map(lamdaA => P(8)(970),lamdaB => P(8)(974),lamdaOut => P(7)(970));
U_F8971: entity F port map(lamdaA => P(8)(971),lamdaB => P(8)(975),lamdaOut => P(7)(971));
U_G8972: entity G port map(lamdaA => P(8)(968),lamdaB => P(8)(972),s => s(8)(484),lamdaOut => P(7)(972));
U_G8973: entity G port map(lamdaA => P(8)(969),lamdaB => P(8)(973),s => s(8)(485),lamdaOut => P(7)(973));
U_G8974: entity G port map(lamdaA => P(8)(970),lamdaB => P(8)(974),s => s(8)(486),lamdaOut => P(7)(974));
U_G8975: entity G port map(lamdaA => P(8)(971),lamdaB => P(8)(975),s => s(8)(487),lamdaOut => P(7)(975));
U_F8976: entity F port map(lamdaA => P(8)(976),lamdaB => P(8)(980),lamdaOut => P(7)(976));
U_F8977: entity F port map(lamdaA => P(8)(977),lamdaB => P(8)(981),lamdaOut => P(7)(977));
U_F8978: entity F port map(lamdaA => P(8)(978),lamdaB => P(8)(982),lamdaOut => P(7)(978));
U_F8979: entity F port map(lamdaA => P(8)(979),lamdaB => P(8)(983),lamdaOut => P(7)(979));
U_G8980: entity G port map(lamdaA => P(8)(976),lamdaB => P(8)(980),s => s(8)(488),lamdaOut => P(7)(980));
U_G8981: entity G port map(lamdaA => P(8)(977),lamdaB => P(8)(981),s => s(8)(489),lamdaOut => P(7)(981));
U_G8982: entity G port map(lamdaA => P(8)(978),lamdaB => P(8)(982),s => s(8)(490),lamdaOut => P(7)(982));
U_G8983: entity G port map(lamdaA => P(8)(979),lamdaB => P(8)(983),s => s(8)(491),lamdaOut => P(7)(983));
U_F8984: entity F port map(lamdaA => P(8)(984),lamdaB => P(8)(988),lamdaOut => P(7)(984));
U_F8985: entity F port map(lamdaA => P(8)(985),lamdaB => P(8)(989),lamdaOut => P(7)(985));
U_F8986: entity F port map(lamdaA => P(8)(986),lamdaB => P(8)(990),lamdaOut => P(7)(986));
U_F8987: entity F port map(lamdaA => P(8)(987),lamdaB => P(8)(991),lamdaOut => P(7)(987));
U_G8988: entity G port map(lamdaA => P(8)(984),lamdaB => P(8)(988),s => s(8)(492),lamdaOut => P(7)(988));
U_G8989: entity G port map(lamdaA => P(8)(985),lamdaB => P(8)(989),s => s(8)(493),lamdaOut => P(7)(989));
U_G8990: entity G port map(lamdaA => P(8)(986),lamdaB => P(8)(990),s => s(8)(494),lamdaOut => P(7)(990));
U_G8991: entity G port map(lamdaA => P(8)(987),lamdaB => P(8)(991),s => s(8)(495),lamdaOut => P(7)(991));
U_F8992: entity F port map(lamdaA => P(8)(992),lamdaB => P(8)(996),lamdaOut => P(7)(992));
U_F8993: entity F port map(lamdaA => P(8)(993),lamdaB => P(8)(997),lamdaOut => P(7)(993));
U_F8994: entity F port map(lamdaA => P(8)(994),lamdaB => P(8)(998),lamdaOut => P(7)(994));
U_F8995: entity F port map(lamdaA => P(8)(995),lamdaB => P(8)(999),lamdaOut => P(7)(995));
U_G8996: entity G port map(lamdaA => P(8)(992),lamdaB => P(8)(996),s => s(8)(496),lamdaOut => P(7)(996));
U_G8997: entity G port map(lamdaA => P(8)(993),lamdaB => P(8)(997),s => s(8)(497),lamdaOut => P(7)(997));
U_G8998: entity G port map(lamdaA => P(8)(994),lamdaB => P(8)(998),s => s(8)(498),lamdaOut => P(7)(998));
U_G8999: entity G port map(lamdaA => P(8)(995),lamdaB => P(8)(999),s => s(8)(499),lamdaOut => P(7)(999));
U_F81000: entity F port map(lamdaA => P(8)(1000),lamdaB => P(8)(1004),lamdaOut => P(7)(1000));
U_F81001: entity F port map(lamdaA => P(8)(1001),lamdaB => P(8)(1005),lamdaOut => P(7)(1001));
U_F81002: entity F port map(lamdaA => P(8)(1002),lamdaB => P(8)(1006),lamdaOut => P(7)(1002));
U_F81003: entity F port map(lamdaA => P(8)(1003),lamdaB => P(8)(1007),lamdaOut => P(7)(1003));
U_G81004: entity G port map(lamdaA => P(8)(1000),lamdaB => P(8)(1004),s => s(8)(500),lamdaOut => P(7)(1004));
U_G81005: entity G port map(lamdaA => P(8)(1001),lamdaB => P(8)(1005),s => s(8)(501),lamdaOut => P(7)(1005));
U_G81006: entity G port map(lamdaA => P(8)(1002),lamdaB => P(8)(1006),s => s(8)(502),lamdaOut => P(7)(1006));
U_G81007: entity G port map(lamdaA => P(8)(1003),lamdaB => P(8)(1007),s => s(8)(503),lamdaOut => P(7)(1007));
U_F81008: entity F port map(lamdaA => P(8)(1008),lamdaB => P(8)(1012),lamdaOut => P(7)(1008));
U_F81009: entity F port map(lamdaA => P(8)(1009),lamdaB => P(8)(1013),lamdaOut => P(7)(1009));
U_F81010: entity F port map(lamdaA => P(8)(1010),lamdaB => P(8)(1014),lamdaOut => P(7)(1010));
U_F81011: entity F port map(lamdaA => P(8)(1011),lamdaB => P(8)(1015),lamdaOut => P(7)(1011));
U_G81012: entity G port map(lamdaA => P(8)(1008),lamdaB => P(8)(1012),s => s(8)(504),lamdaOut => P(7)(1012));
U_G81013: entity G port map(lamdaA => P(8)(1009),lamdaB => P(8)(1013),s => s(8)(505),lamdaOut => P(7)(1013));
U_G81014: entity G port map(lamdaA => P(8)(1010),lamdaB => P(8)(1014),s => s(8)(506),lamdaOut => P(7)(1014));
U_G81015: entity G port map(lamdaA => P(8)(1011),lamdaB => P(8)(1015),s => s(8)(507),lamdaOut => P(7)(1015));
U_F81016: entity F port map(lamdaA => P(8)(1016),lamdaB => P(8)(1020),lamdaOut => P(7)(1016));
U_F81017: entity F port map(lamdaA => P(8)(1017),lamdaB => P(8)(1021),lamdaOut => P(7)(1017));
U_F81018: entity F port map(lamdaA => P(8)(1018),lamdaB => P(8)(1022),lamdaOut => P(7)(1018));
U_F81019: entity F port map(lamdaA => P(8)(1019),lamdaB => P(8)(1023),lamdaOut => P(7)(1019));
U_G81020: entity G port map(lamdaA => P(8)(1016),lamdaB => P(8)(1020),s => s(8)(508),lamdaOut => P(7)(1020));
U_G81021: entity G port map(lamdaA => P(8)(1017),lamdaB => P(8)(1021),s => s(8)(509),lamdaOut => P(7)(1021));
U_G81022: entity G port map(lamdaA => P(8)(1018),lamdaB => P(8)(1022),s => s(8)(510),lamdaOut => P(7)(1022));
U_G81023: entity G port map(lamdaA => P(8)(1019),lamdaB => P(8)(1023),s => s(8)(511),lamdaOut => P(7)(1023));
-- STAGE 6
U_F70: entity F port map(lamdaA => P(7)(0),lamdaB => P(7)(8),lamdaOut => P(6)(0));
U_F71: entity F port map(lamdaA => P(7)(1),lamdaB => P(7)(9),lamdaOut => P(6)(1));
U_F72: entity F port map(lamdaA => P(7)(2),lamdaB => P(7)(10),lamdaOut => P(6)(2));
U_F73: entity F port map(lamdaA => P(7)(3),lamdaB => P(7)(11),lamdaOut => P(6)(3));
U_F74: entity F port map(lamdaA => P(7)(4),lamdaB => P(7)(12),lamdaOut => P(6)(4));
U_F75: entity F port map(lamdaA => P(7)(5),lamdaB => P(7)(13),lamdaOut => P(6)(5));
U_F76: entity F port map(lamdaA => P(7)(6),lamdaB => P(7)(14),lamdaOut => P(6)(6));
U_F77: entity F port map(lamdaA => P(7)(7),lamdaB => P(7)(15),lamdaOut => P(6)(7));
U_G78: entity G port map(lamdaA => P(7)(0),lamdaB => P(7)(8),s => s(7)(0),lamdaOut => P(6)(8));
U_G79: entity G port map(lamdaA => P(7)(1),lamdaB => P(7)(9),s => s(7)(1),lamdaOut => P(6)(9));
U_G710: entity G port map(lamdaA => P(7)(2),lamdaB => P(7)(10),s => s(7)(2),lamdaOut => P(6)(10));
U_G711: entity G port map(lamdaA => P(7)(3),lamdaB => P(7)(11),s => s(7)(3),lamdaOut => P(6)(11));
U_G712: entity G port map(lamdaA => P(7)(4),lamdaB => P(7)(12),s => s(7)(4),lamdaOut => P(6)(12));
U_G713: entity G port map(lamdaA => P(7)(5),lamdaB => P(7)(13),s => s(7)(5),lamdaOut => P(6)(13));
U_G714: entity G port map(lamdaA => P(7)(6),lamdaB => P(7)(14),s => s(7)(6),lamdaOut => P(6)(14));
U_G715: entity G port map(lamdaA => P(7)(7),lamdaB => P(7)(15),s => s(7)(7),lamdaOut => P(6)(15));
U_F716: entity F port map(lamdaA => P(7)(16),lamdaB => P(7)(24),lamdaOut => P(6)(16));
U_F717: entity F port map(lamdaA => P(7)(17),lamdaB => P(7)(25),lamdaOut => P(6)(17));
U_F718: entity F port map(lamdaA => P(7)(18),lamdaB => P(7)(26),lamdaOut => P(6)(18));
U_F719: entity F port map(lamdaA => P(7)(19),lamdaB => P(7)(27),lamdaOut => P(6)(19));
U_F720: entity F port map(lamdaA => P(7)(20),lamdaB => P(7)(28),lamdaOut => P(6)(20));
U_F721: entity F port map(lamdaA => P(7)(21),lamdaB => P(7)(29),lamdaOut => P(6)(21));
U_F722: entity F port map(lamdaA => P(7)(22),lamdaB => P(7)(30),lamdaOut => P(6)(22));
U_F723: entity F port map(lamdaA => P(7)(23),lamdaB => P(7)(31),lamdaOut => P(6)(23));
U_G724: entity G port map(lamdaA => P(7)(16),lamdaB => P(7)(24),s => s(7)(8),lamdaOut => P(6)(24));
U_G725: entity G port map(lamdaA => P(7)(17),lamdaB => P(7)(25),s => s(7)(9),lamdaOut => P(6)(25));
U_G726: entity G port map(lamdaA => P(7)(18),lamdaB => P(7)(26),s => s(7)(10),lamdaOut => P(6)(26));
U_G727: entity G port map(lamdaA => P(7)(19),lamdaB => P(7)(27),s => s(7)(11),lamdaOut => P(6)(27));
U_G728: entity G port map(lamdaA => P(7)(20),lamdaB => P(7)(28),s => s(7)(12),lamdaOut => P(6)(28));
U_G729: entity G port map(lamdaA => P(7)(21),lamdaB => P(7)(29),s => s(7)(13),lamdaOut => P(6)(29));
U_G730: entity G port map(lamdaA => P(7)(22),lamdaB => P(7)(30),s => s(7)(14),lamdaOut => P(6)(30));
U_G731: entity G port map(lamdaA => P(7)(23),lamdaB => P(7)(31),s => s(7)(15),lamdaOut => P(6)(31));
U_F732: entity F port map(lamdaA => P(7)(32),lamdaB => P(7)(40),lamdaOut => P(6)(32));
U_F733: entity F port map(lamdaA => P(7)(33),lamdaB => P(7)(41),lamdaOut => P(6)(33));
U_F734: entity F port map(lamdaA => P(7)(34),lamdaB => P(7)(42),lamdaOut => P(6)(34));
U_F735: entity F port map(lamdaA => P(7)(35),lamdaB => P(7)(43),lamdaOut => P(6)(35));
U_F736: entity F port map(lamdaA => P(7)(36),lamdaB => P(7)(44),lamdaOut => P(6)(36));
U_F737: entity F port map(lamdaA => P(7)(37),lamdaB => P(7)(45),lamdaOut => P(6)(37));
U_F738: entity F port map(lamdaA => P(7)(38),lamdaB => P(7)(46),lamdaOut => P(6)(38));
U_F739: entity F port map(lamdaA => P(7)(39),lamdaB => P(7)(47),lamdaOut => P(6)(39));
U_G740: entity G port map(lamdaA => P(7)(32),lamdaB => P(7)(40),s => s(7)(16),lamdaOut => P(6)(40));
U_G741: entity G port map(lamdaA => P(7)(33),lamdaB => P(7)(41),s => s(7)(17),lamdaOut => P(6)(41));
U_G742: entity G port map(lamdaA => P(7)(34),lamdaB => P(7)(42),s => s(7)(18),lamdaOut => P(6)(42));
U_G743: entity G port map(lamdaA => P(7)(35),lamdaB => P(7)(43),s => s(7)(19),lamdaOut => P(6)(43));
U_G744: entity G port map(lamdaA => P(7)(36),lamdaB => P(7)(44),s => s(7)(20),lamdaOut => P(6)(44));
U_G745: entity G port map(lamdaA => P(7)(37),lamdaB => P(7)(45),s => s(7)(21),lamdaOut => P(6)(45));
U_G746: entity G port map(lamdaA => P(7)(38),lamdaB => P(7)(46),s => s(7)(22),lamdaOut => P(6)(46));
U_G747: entity G port map(lamdaA => P(7)(39),lamdaB => P(7)(47),s => s(7)(23),lamdaOut => P(6)(47));
U_F748: entity F port map(lamdaA => P(7)(48),lamdaB => P(7)(56),lamdaOut => P(6)(48));
U_F749: entity F port map(lamdaA => P(7)(49),lamdaB => P(7)(57),lamdaOut => P(6)(49));
U_F750: entity F port map(lamdaA => P(7)(50),lamdaB => P(7)(58),lamdaOut => P(6)(50));
U_F751: entity F port map(lamdaA => P(7)(51),lamdaB => P(7)(59),lamdaOut => P(6)(51));
U_F752: entity F port map(lamdaA => P(7)(52),lamdaB => P(7)(60),lamdaOut => P(6)(52));
U_F753: entity F port map(lamdaA => P(7)(53),lamdaB => P(7)(61),lamdaOut => P(6)(53));
U_F754: entity F port map(lamdaA => P(7)(54),lamdaB => P(7)(62),lamdaOut => P(6)(54));
U_F755: entity F port map(lamdaA => P(7)(55),lamdaB => P(7)(63),lamdaOut => P(6)(55));
U_G756: entity G port map(lamdaA => P(7)(48),lamdaB => P(7)(56),s => s(7)(24),lamdaOut => P(6)(56));
U_G757: entity G port map(lamdaA => P(7)(49),lamdaB => P(7)(57),s => s(7)(25),lamdaOut => P(6)(57));
U_G758: entity G port map(lamdaA => P(7)(50),lamdaB => P(7)(58),s => s(7)(26),lamdaOut => P(6)(58));
U_G759: entity G port map(lamdaA => P(7)(51),lamdaB => P(7)(59),s => s(7)(27),lamdaOut => P(6)(59));
U_G760: entity G port map(lamdaA => P(7)(52),lamdaB => P(7)(60),s => s(7)(28),lamdaOut => P(6)(60));
U_G761: entity G port map(lamdaA => P(7)(53),lamdaB => P(7)(61),s => s(7)(29),lamdaOut => P(6)(61));
U_G762: entity G port map(lamdaA => P(7)(54),lamdaB => P(7)(62),s => s(7)(30),lamdaOut => P(6)(62));
U_G763: entity G port map(lamdaA => P(7)(55),lamdaB => P(7)(63),s => s(7)(31),lamdaOut => P(6)(63));
U_F764: entity F port map(lamdaA => P(7)(64),lamdaB => P(7)(72),lamdaOut => P(6)(64));
U_F765: entity F port map(lamdaA => P(7)(65),lamdaB => P(7)(73),lamdaOut => P(6)(65));
U_F766: entity F port map(lamdaA => P(7)(66),lamdaB => P(7)(74),lamdaOut => P(6)(66));
U_F767: entity F port map(lamdaA => P(7)(67),lamdaB => P(7)(75),lamdaOut => P(6)(67));
U_F768: entity F port map(lamdaA => P(7)(68),lamdaB => P(7)(76),lamdaOut => P(6)(68));
U_F769: entity F port map(lamdaA => P(7)(69),lamdaB => P(7)(77),lamdaOut => P(6)(69));
U_F770: entity F port map(lamdaA => P(7)(70),lamdaB => P(7)(78),lamdaOut => P(6)(70));
U_F771: entity F port map(lamdaA => P(7)(71),lamdaB => P(7)(79),lamdaOut => P(6)(71));
U_G772: entity G port map(lamdaA => P(7)(64),lamdaB => P(7)(72),s => s(7)(32),lamdaOut => P(6)(72));
U_G773: entity G port map(lamdaA => P(7)(65),lamdaB => P(7)(73),s => s(7)(33),lamdaOut => P(6)(73));
U_G774: entity G port map(lamdaA => P(7)(66),lamdaB => P(7)(74),s => s(7)(34),lamdaOut => P(6)(74));
U_G775: entity G port map(lamdaA => P(7)(67),lamdaB => P(7)(75),s => s(7)(35),lamdaOut => P(6)(75));
U_G776: entity G port map(lamdaA => P(7)(68),lamdaB => P(7)(76),s => s(7)(36),lamdaOut => P(6)(76));
U_G777: entity G port map(lamdaA => P(7)(69),lamdaB => P(7)(77),s => s(7)(37),lamdaOut => P(6)(77));
U_G778: entity G port map(lamdaA => P(7)(70),lamdaB => P(7)(78),s => s(7)(38),lamdaOut => P(6)(78));
U_G779: entity G port map(lamdaA => P(7)(71),lamdaB => P(7)(79),s => s(7)(39),lamdaOut => P(6)(79));
U_F780: entity F port map(lamdaA => P(7)(80),lamdaB => P(7)(88),lamdaOut => P(6)(80));
U_F781: entity F port map(lamdaA => P(7)(81),lamdaB => P(7)(89),lamdaOut => P(6)(81));
U_F782: entity F port map(lamdaA => P(7)(82),lamdaB => P(7)(90),lamdaOut => P(6)(82));
U_F783: entity F port map(lamdaA => P(7)(83),lamdaB => P(7)(91),lamdaOut => P(6)(83));
U_F784: entity F port map(lamdaA => P(7)(84),lamdaB => P(7)(92),lamdaOut => P(6)(84));
U_F785: entity F port map(lamdaA => P(7)(85),lamdaB => P(7)(93),lamdaOut => P(6)(85));
U_F786: entity F port map(lamdaA => P(7)(86),lamdaB => P(7)(94),lamdaOut => P(6)(86));
U_F787: entity F port map(lamdaA => P(7)(87),lamdaB => P(7)(95),lamdaOut => P(6)(87));
U_G788: entity G port map(lamdaA => P(7)(80),lamdaB => P(7)(88),s => s(7)(40),lamdaOut => P(6)(88));
U_G789: entity G port map(lamdaA => P(7)(81),lamdaB => P(7)(89),s => s(7)(41),lamdaOut => P(6)(89));
U_G790: entity G port map(lamdaA => P(7)(82),lamdaB => P(7)(90),s => s(7)(42),lamdaOut => P(6)(90));
U_G791: entity G port map(lamdaA => P(7)(83),lamdaB => P(7)(91),s => s(7)(43),lamdaOut => P(6)(91));
U_G792: entity G port map(lamdaA => P(7)(84),lamdaB => P(7)(92),s => s(7)(44),lamdaOut => P(6)(92));
U_G793: entity G port map(lamdaA => P(7)(85),lamdaB => P(7)(93),s => s(7)(45),lamdaOut => P(6)(93));
U_G794: entity G port map(lamdaA => P(7)(86),lamdaB => P(7)(94),s => s(7)(46),lamdaOut => P(6)(94));
U_G795: entity G port map(lamdaA => P(7)(87),lamdaB => P(7)(95),s => s(7)(47),lamdaOut => P(6)(95));
U_F796: entity F port map(lamdaA => P(7)(96),lamdaB => P(7)(104),lamdaOut => P(6)(96));
U_F797: entity F port map(lamdaA => P(7)(97),lamdaB => P(7)(105),lamdaOut => P(6)(97));
U_F798: entity F port map(lamdaA => P(7)(98),lamdaB => P(7)(106),lamdaOut => P(6)(98));
U_F799: entity F port map(lamdaA => P(7)(99),lamdaB => P(7)(107),lamdaOut => P(6)(99));
U_F7100: entity F port map(lamdaA => P(7)(100),lamdaB => P(7)(108),lamdaOut => P(6)(100));
U_F7101: entity F port map(lamdaA => P(7)(101),lamdaB => P(7)(109),lamdaOut => P(6)(101));
U_F7102: entity F port map(lamdaA => P(7)(102),lamdaB => P(7)(110),lamdaOut => P(6)(102));
U_F7103: entity F port map(lamdaA => P(7)(103),lamdaB => P(7)(111),lamdaOut => P(6)(103));
U_G7104: entity G port map(lamdaA => P(7)(96),lamdaB => P(7)(104),s => s(7)(48),lamdaOut => P(6)(104));
U_G7105: entity G port map(lamdaA => P(7)(97),lamdaB => P(7)(105),s => s(7)(49),lamdaOut => P(6)(105));
U_G7106: entity G port map(lamdaA => P(7)(98),lamdaB => P(7)(106),s => s(7)(50),lamdaOut => P(6)(106));
U_G7107: entity G port map(lamdaA => P(7)(99),lamdaB => P(7)(107),s => s(7)(51),lamdaOut => P(6)(107));
U_G7108: entity G port map(lamdaA => P(7)(100),lamdaB => P(7)(108),s => s(7)(52),lamdaOut => P(6)(108));
U_G7109: entity G port map(lamdaA => P(7)(101),lamdaB => P(7)(109),s => s(7)(53),lamdaOut => P(6)(109));
U_G7110: entity G port map(lamdaA => P(7)(102),lamdaB => P(7)(110),s => s(7)(54),lamdaOut => P(6)(110));
U_G7111: entity G port map(lamdaA => P(7)(103),lamdaB => P(7)(111),s => s(7)(55),lamdaOut => P(6)(111));
U_F7112: entity F port map(lamdaA => P(7)(112),lamdaB => P(7)(120),lamdaOut => P(6)(112));
U_F7113: entity F port map(lamdaA => P(7)(113),lamdaB => P(7)(121),lamdaOut => P(6)(113));
U_F7114: entity F port map(lamdaA => P(7)(114),lamdaB => P(7)(122),lamdaOut => P(6)(114));
U_F7115: entity F port map(lamdaA => P(7)(115),lamdaB => P(7)(123),lamdaOut => P(6)(115));
U_F7116: entity F port map(lamdaA => P(7)(116),lamdaB => P(7)(124),lamdaOut => P(6)(116));
U_F7117: entity F port map(lamdaA => P(7)(117),lamdaB => P(7)(125),lamdaOut => P(6)(117));
U_F7118: entity F port map(lamdaA => P(7)(118),lamdaB => P(7)(126),lamdaOut => P(6)(118));
U_F7119: entity F port map(lamdaA => P(7)(119),lamdaB => P(7)(127),lamdaOut => P(6)(119));
U_G7120: entity G port map(lamdaA => P(7)(112),lamdaB => P(7)(120),s => s(7)(56),lamdaOut => P(6)(120));
U_G7121: entity G port map(lamdaA => P(7)(113),lamdaB => P(7)(121),s => s(7)(57),lamdaOut => P(6)(121));
U_G7122: entity G port map(lamdaA => P(7)(114),lamdaB => P(7)(122),s => s(7)(58),lamdaOut => P(6)(122));
U_G7123: entity G port map(lamdaA => P(7)(115),lamdaB => P(7)(123),s => s(7)(59),lamdaOut => P(6)(123));
U_G7124: entity G port map(lamdaA => P(7)(116),lamdaB => P(7)(124),s => s(7)(60),lamdaOut => P(6)(124));
U_G7125: entity G port map(lamdaA => P(7)(117),lamdaB => P(7)(125),s => s(7)(61),lamdaOut => P(6)(125));
U_G7126: entity G port map(lamdaA => P(7)(118),lamdaB => P(7)(126),s => s(7)(62),lamdaOut => P(6)(126));
U_G7127: entity G port map(lamdaA => P(7)(119),lamdaB => P(7)(127),s => s(7)(63),lamdaOut => P(6)(127));
U_F7128: entity F port map(lamdaA => P(7)(128),lamdaB => P(7)(136),lamdaOut => P(6)(128));
U_F7129: entity F port map(lamdaA => P(7)(129),lamdaB => P(7)(137),lamdaOut => P(6)(129));
U_F7130: entity F port map(lamdaA => P(7)(130),lamdaB => P(7)(138),lamdaOut => P(6)(130));
U_F7131: entity F port map(lamdaA => P(7)(131),lamdaB => P(7)(139),lamdaOut => P(6)(131));
U_F7132: entity F port map(lamdaA => P(7)(132),lamdaB => P(7)(140),lamdaOut => P(6)(132));
U_F7133: entity F port map(lamdaA => P(7)(133),lamdaB => P(7)(141),lamdaOut => P(6)(133));
U_F7134: entity F port map(lamdaA => P(7)(134),lamdaB => P(7)(142),lamdaOut => P(6)(134));
U_F7135: entity F port map(lamdaA => P(7)(135),lamdaB => P(7)(143),lamdaOut => P(6)(135));
U_G7136: entity G port map(lamdaA => P(7)(128),lamdaB => P(7)(136),s => s(7)(64),lamdaOut => P(6)(136));
U_G7137: entity G port map(lamdaA => P(7)(129),lamdaB => P(7)(137),s => s(7)(65),lamdaOut => P(6)(137));
U_G7138: entity G port map(lamdaA => P(7)(130),lamdaB => P(7)(138),s => s(7)(66),lamdaOut => P(6)(138));
U_G7139: entity G port map(lamdaA => P(7)(131),lamdaB => P(7)(139),s => s(7)(67),lamdaOut => P(6)(139));
U_G7140: entity G port map(lamdaA => P(7)(132),lamdaB => P(7)(140),s => s(7)(68),lamdaOut => P(6)(140));
U_G7141: entity G port map(lamdaA => P(7)(133),lamdaB => P(7)(141),s => s(7)(69),lamdaOut => P(6)(141));
U_G7142: entity G port map(lamdaA => P(7)(134),lamdaB => P(7)(142),s => s(7)(70),lamdaOut => P(6)(142));
U_G7143: entity G port map(lamdaA => P(7)(135),lamdaB => P(7)(143),s => s(7)(71),lamdaOut => P(6)(143));
U_F7144: entity F port map(lamdaA => P(7)(144),lamdaB => P(7)(152),lamdaOut => P(6)(144));
U_F7145: entity F port map(lamdaA => P(7)(145),lamdaB => P(7)(153),lamdaOut => P(6)(145));
U_F7146: entity F port map(lamdaA => P(7)(146),lamdaB => P(7)(154),lamdaOut => P(6)(146));
U_F7147: entity F port map(lamdaA => P(7)(147),lamdaB => P(7)(155),lamdaOut => P(6)(147));
U_F7148: entity F port map(lamdaA => P(7)(148),lamdaB => P(7)(156),lamdaOut => P(6)(148));
U_F7149: entity F port map(lamdaA => P(7)(149),lamdaB => P(7)(157),lamdaOut => P(6)(149));
U_F7150: entity F port map(lamdaA => P(7)(150),lamdaB => P(7)(158),lamdaOut => P(6)(150));
U_F7151: entity F port map(lamdaA => P(7)(151),lamdaB => P(7)(159),lamdaOut => P(6)(151));
U_G7152: entity G port map(lamdaA => P(7)(144),lamdaB => P(7)(152),s => s(7)(72),lamdaOut => P(6)(152));
U_G7153: entity G port map(lamdaA => P(7)(145),lamdaB => P(7)(153),s => s(7)(73),lamdaOut => P(6)(153));
U_G7154: entity G port map(lamdaA => P(7)(146),lamdaB => P(7)(154),s => s(7)(74),lamdaOut => P(6)(154));
U_G7155: entity G port map(lamdaA => P(7)(147),lamdaB => P(7)(155),s => s(7)(75),lamdaOut => P(6)(155));
U_G7156: entity G port map(lamdaA => P(7)(148),lamdaB => P(7)(156),s => s(7)(76),lamdaOut => P(6)(156));
U_G7157: entity G port map(lamdaA => P(7)(149),lamdaB => P(7)(157),s => s(7)(77),lamdaOut => P(6)(157));
U_G7158: entity G port map(lamdaA => P(7)(150),lamdaB => P(7)(158),s => s(7)(78),lamdaOut => P(6)(158));
U_G7159: entity G port map(lamdaA => P(7)(151),lamdaB => P(7)(159),s => s(7)(79),lamdaOut => P(6)(159));
U_F7160: entity F port map(lamdaA => P(7)(160),lamdaB => P(7)(168),lamdaOut => P(6)(160));
U_F7161: entity F port map(lamdaA => P(7)(161),lamdaB => P(7)(169),lamdaOut => P(6)(161));
U_F7162: entity F port map(lamdaA => P(7)(162),lamdaB => P(7)(170),lamdaOut => P(6)(162));
U_F7163: entity F port map(lamdaA => P(7)(163),lamdaB => P(7)(171),lamdaOut => P(6)(163));
U_F7164: entity F port map(lamdaA => P(7)(164),lamdaB => P(7)(172),lamdaOut => P(6)(164));
U_F7165: entity F port map(lamdaA => P(7)(165),lamdaB => P(7)(173),lamdaOut => P(6)(165));
U_F7166: entity F port map(lamdaA => P(7)(166),lamdaB => P(7)(174),lamdaOut => P(6)(166));
U_F7167: entity F port map(lamdaA => P(7)(167),lamdaB => P(7)(175),lamdaOut => P(6)(167));
U_G7168: entity G port map(lamdaA => P(7)(160),lamdaB => P(7)(168),s => s(7)(80),lamdaOut => P(6)(168));
U_G7169: entity G port map(lamdaA => P(7)(161),lamdaB => P(7)(169),s => s(7)(81),lamdaOut => P(6)(169));
U_G7170: entity G port map(lamdaA => P(7)(162),lamdaB => P(7)(170),s => s(7)(82),lamdaOut => P(6)(170));
U_G7171: entity G port map(lamdaA => P(7)(163),lamdaB => P(7)(171),s => s(7)(83),lamdaOut => P(6)(171));
U_G7172: entity G port map(lamdaA => P(7)(164),lamdaB => P(7)(172),s => s(7)(84),lamdaOut => P(6)(172));
U_G7173: entity G port map(lamdaA => P(7)(165),lamdaB => P(7)(173),s => s(7)(85),lamdaOut => P(6)(173));
U_G7174: entity G port map(lamdaA => P(7)(166),lamdaB => P(7)(174),s => s(7)(86),lamdaOut => P(6)(174));
U_G7175: entity G port map(lamdaA => P(7)(167),lamdaB => P(7)(175),s => s(7)(87),lamdaOut => P(6)(175));
U_F7176: entity F port map(lamdaA => P(7)(176),lamdaB => P(7)(184),lamdaOut => P(6)(176));
U_F7177: entity F port map(lamdaA => P(7)(177),lamdaB => P(7)(185),lamdaOut => P(6)(177));
U_F7178: entity F port map(lamdaA => P(7)(178),lamdaB => P(7)(186),lamdaOut => P(6)(178));
U_F7179: entity F port map(lamdaA => P(7)(179),lamdaB => P(7)(187),lamdaOut => P(6)(179));
U_F7180: entity F port map(lamdaA => P(7)(180),lamdaB => P(7)(188),lamdaOut => P(6)(180));
U_F7181: entity F port map(lamdaA => P(7)(181),lamdaB => P(7)(189),lamdaOut => P(6)(181));
U_F7182: entity F port map(lamdaA => P(7)(182),lamdaB => P(7)(190),lamdaOut => P(6)(182));
U_F7183: entity F port map(lamdaA => P(7)(183),lamdaB => P(7)(191),lamdaOut => P(6)(183));
U_G7184: entity G port map(lamdaA => P(7)(176),lamdaB => P(7)(184),s => s(7)(88),lamdaOut => P(6)(184));
U_G7185: entity G port map(lamdaA => P(7)(177),lamdaB => P(7)(185),s => s(7)(89),lamdaOut => P(6)(185));
U_G7186: entity G port map(lamdaA => P(7)(178),lamdaB => P(7)(186),s => s(7)(90),lamdaOut => P(6)(186));
U_G7187: entity G port map(lamdaA => P(7)(179),lamdaB => P(7)(187),s => s(7)(91),lamdaOut => P(6)(187));
U_G7188: entity G port map(lamdaA => P(7)(180),lamdaB => P(7)(188),s => s(7)(92),lamdaOut => P(6)(188));
U_G7189: entity G port map(lamdaA => P(7)(181),lamdaB => P(7)(189),s => s(7)(93),lamdaOut => P(6)(189));
U_G7190: entity G port map(lamdaA => P(7)(182),lamdaB => P(7)(190),s => s(7)(94),lamdaOut => P(6)(190));
U_G7191: entity G port map(lamdaA => P(7)(183),lamdaB => P(7)(191),s => s(7)(95),lamdaOut => P(6)(191));
U_F7192: entity F port map(lamdaA => P(7)(192),lamdaB => P(7)(200),lamdaOut => P(6)(192));
U_F7193: entity F port map(lamdaA => P(7)(193),lamdaB => P(7)(201),lamdaOut => P(6)(193));
U_F7194: entity F port map(lamdaA => P(7)(194),lamdaB => P(7)(202),lamdaOut => P(6)(194));
U_F7195: entity F port map(lamdaA => P(7)(195),lamdaB => P(7)(203),lamdaOut => P(6)(195));
U_F7196: entity F port map(lamdaA => P(7)(196),lamdaB => P(7)(204),lamdaOut => P(6)(196));
U_F7197: entity F port map(lamdaA => P(7)(197),lamdaB => P(7)(205),lamdaOut => P(6)(197));
U_F7198: entity F port map(lamdaA => P(7)(198),lamdaB => P(7)(206),lamdaOut => P(6)(198));
U_F7199: entity F port map(lamdaA => P(7)(199),lamdaB => P(7)(207),lamdaOut => P(6)(199));
U_G7200: entity G port map(lamdaA => P(7)(192),lamdaB => P(7)(200),s => s(7)(96),lamdaOut => P(6)(200));
U_G7201: entity G port map(lamdaA => P(7)(193),lamdaB => P(7)(201),s => s(7)(97),lamdaOut => P(6)(201));
U_G7202: entity G port map(lamdaA => P(7)(194),lamdaB => P(7)(202),s => s(7)(98),lamdaOut => P(6)(202));
U_G7203: entity G port map(lamdaA => P(7)(195),lamdaB => P(7)(203),s => s(7)(99),lamdaOut => P(6)(203));
U_G7204: entity G port map(lamdaA => P(7)(196),lamdaB => P(7)(204),s => s(7)(100),lamdaOut => P(6)(204));
U_G7205: entity G port map(lamdaA => P(7)(197),lamdaB => P(7)(205),s => s(7)(101),lamdaOut => P(6)(205));
U_G7206: entity G port map(lamdaA => P(7)(198),lamdaB => P(7)(206),s => s(7)(102),lamdaOut => P(6)(206));
U_G7207: entity G port map(lamdaA => P(7)(199),lamdaB => P(7)(207),s => s(7)(103),lamdaOut => P(6)(207));
U_F7208: entity F port map(lamdaA => P(7)(208),lamdaB => P(7)(216),lamdaOut => P(6)(208));
U_F7209: entity F port map(lamdaA => P(7)(209),lamdaB => P(7)(217),lamdaOut => P(6)(209));
U_F7210: entity F port map(lamdaA => P(7)(210),lamdaB => P(7)(218),lamdaOut => P(6)(210));
U_F7211: entity F port map(lamdaA => P(7)(211),lamdaB => P(7)(219),lamdaOut => P(6)(211));
U_F7212: entity F port map(lamdaA => P(7)(212),lamdaB => P(7)(220),lamdaOut => P(6)(212));
U_F7213: entity F port map(lamdaA => P(7)(213),lamdaB => P(7)(221),lamdaOut => P(6)(213));
U_F7214: entity F port map(lamdaA => P(7)(214),lamdaB => P(7)(222),lamdaOut => P(6)(214));
U_F7215: entity F port map(lamdaA => P(7)(215),lamdaB => P(7)(223),lamdaOut => P(6)(215));
U_G7216: entity G port map(lamdaA => P(7)(208),lamdaB => P(7)(216),s => s(7)(104),lamdaOut => P(6)(216));
U_G7217: entity G port map(lamdaA => P(7)(209),lamdaB => P(7)(217),s => s(7)(105),lamdaOut => P(6)(217));
U_G7218: entity G port map(lamdaA => P(7)(210),lamdaB => P(7)(218),s => s(7)(106),lamdaOut => P(6)(218));
U_G7219: entity G port map(lamdaA => P(7)(211),lamdaB => P(7)(219),s => s(7)(107),lamdaOut => P(6)(219));
U_G7220: entity G port map(lamdaA => P(7)(212),lamdaB => P(7)(220),s => s(7)(108),lamdaOut => P(6)(220));
U_G7221: entity G port map(lamdaA => P(7)(213),lamdaB => P(7)(221),s => s(7)(109),lamdaOut => P(6)(221));
U_G7222: entity G port map(lamdaA => P(7)(214),lamdaB => P(7)(222),s => s(7)(110),lamdaOut => P(6)(222));
U_G7223: entity G port map(lamdaA => P(7)(215),lamdaB => P(7)(223),s => s(7)(111),lamdaOut => P(6)(223));
U_F7224: entity F port map(lamdaA => P(7)(224),lamdaB => P(7)(232),lamdaOut => P(6)(224));
U_F7225: entity F port map(lamdaA => P(7)(225),lamdaB => P(7)(233),lamdaOut => P(6)(225));
U_F7226: entity F port map(lamdaA => P(7)(226),lamdaB => P(7)(234),lamdaOut => P(6)(226));
U_F7227: entity F port map(lamdaA => P(7)(227),lamdaB => P(7)(235),lamdaOut => P(6)(227));
U_F7228: entity F port map(lamdaA => P(7)(228),lamdaB => P(7)(236),lamdaOut => P(6)(228));
U_F7229: entity F port map(lamdaA => P(7)(229),lamdaB => P(7)(237),lamdaOut => P(6)(229));
U_F7230: entity F port map(lamdaA => P(7)(230),lamdaB => P(7)(238),lamdaOut => P(6)(230));
U_F7231: entity F port map(lamdaA => P(7)(231),lamdaB => P(7)(239),lamdaOut => P(6)(231));
U_G7232: entity G port map(lamdaA => P(7)(224),lamdaB => P(7)(232),s => s(7)(112),lamdaOut => P(6)(232));
U_G7233: entity G port map(lamdaA => P(7)(225),lamdaB => P(7)(233),s => s(7)(113),lamdaOut => P(6)(233));
U_G7234: entity G port map(lamdaA => P(7)(226),lamdaB => P(7)(234),s => s(7)(114),lamdaOut => P(6)(234));
U_G7235: entity G port map(lamdaA => P(7)(227),lamdaB => P(7)(235),s => s(7)(115),lamdaOut => P(6)(235));
U_G7236: entity G port map(lamdaA => P(7)(228),lamdaB => P(7)(236),s => s(7)(116),lamdaOut => P(6)(236));
U_G7237: entity G port map(lamdaA => P(7)(229),lamdaB => P(7)(237),s => s(7)(117),lamdaOut => P(6)(237));
U_G7238: entity G port map(lamdaA => P(7)(230),lamdaB => P(7)(238),s => s(7)(118),lamdaOut => P(6)(238));
U_G7239: entity G port map(lamdaA => P(7)(231),lamdaB => P(7)(239),s => s(7)(119),lamdaOut => P(6)(239));
U_F7240: entity F port map(lamdaA => P(7)(240),lamdaB => P(7)(248),lamdaOut => P(6)(240));
U_F7241: entity F port map(lamdaA => P(7)(241),lamdaB => P(7)(249),lamdaOut => P(6)(241));
U_F7242: entity F port map(lamdaA => P(7)(242),lamdaB => P(7)(250),lamdaOut => P(6)(242));
U_F7243: entity F port map(lamdaA => P(7)(243),lamdaB => P(7)(251),lamdaOut => P(6)(243));
U_F7244: entity F port map(lamdaA => P(7)(244),lamdaB => P(7)(252),lamdaOut => P(6)(244));
U_F7245: entity F port map(lamdaA => P(7)(245),lamdaB => P(7)(253),lamdaOut => P(6)(245));
U_F7246: entity F port map(lamdaA => P(7)(246),lamdaB => P(7)(254),lamdaOut => P(6)(246));
U_F7247: entity F port map(lamdaA => P(7)(247),lamdaB => P(7)(255),lamdaOut => P(6)(247));
U_G7248: entity G port map(lamdaA => P(7)(240),lamdaB => P(7)(248),s => s(7)(120),lamdaOut => P(6)(248));
U_G7249: entity G port map(lamdaA => P(7)(241),lamdaB => P(7)(249),s => s(7)(121),lamdaOut => P(6)(249));
U_G7250: entity G port map(lamdaA => P(7)(242),lamdaB => P(7)(250),s => s(7)(122),lamdaOut => P(6)(250));
U_G7251: entity G port map(lamdaA => P(7)(243),lamdaB => P(7)(251),s => s(7)(123),lamdaOut => P(6)(251));
U_G7252: entity G port map(lamdaA => P(7)(244),lamdaB => P(7)(252),s => s(7)(124),lamdaOut => P(6)(252));
U_G7253: entity G port map(lamdaA => P(7)(245),lamdaB => P(7)(253),s => s(7)(125),lamdaOut => P(6)(253));
U_G7254: entity G port map(lamdaA => P(7)(246),lamdaB => P(7)(254),s => s(7)(126),lamdaOut => P(6)(254));
U_G7255: entity G port map(lamdaA => P(7)(247),lamdaB => P(7)(255),s => s(7)(127),lamdaOut => P(6)(255));
U_F7256: entity F port map(lamdaA => P(7)(256),lamdaB => P(7)(264),lamdaOut => P(6)(256));
U_F7257: entity F port map(lamdaA => P(7)(257),lamdaB => P(7)(265),lamdaOut => P(6)(257));
U_F7258: entity F port map(lamdaA => P(7)(258),lamdaB => P(7)(266),lamdaOut => P(6)(258));
U_F7259: entity F port map(lamdaA => P(7)(259),lamdaB => P(7)(267),lamdaOut => P(6)(259));
U_F7260: entity F port map(lamdaA => P(7)(260),lamdaB => P(7)(268),lamdaOut => P(6)(260));
U_F7261: entity F port map(lamdaA => P(7)(261),lamdaB => P(7)(269),lamdaOut => P(6)(261));
U_F7262: entity F port map(lamdaA => P(7)(262),lamdaB => P(7)(270),lamdaOut => P(6)(262));
U_F7263: entity F port map(lamdaA => P(7)(263),lamdaB => P(7)(271),lamdaOut => P(6)(263));
U_G7264: entity G port map(lamdaA => P(7)(256),lamdaB => P(7)(264),s => s(7)(128),lamdaOut => P(6)(264));
U_G7265: entity G port map(lamdaA => P(7)(257),lamdaB => P(7)(265),s => s(7)(129),lamdaOut => P(6)(265));
U_G7266: entity G port map(lamdaA => P(7)(258),lamdaB => P(7)(266),s => s(7)(130),lamdaOut => P(6)(266));
U_G7267: entity G port map(lamdaA => P(7)(259),lamdaB => P(7)(267),s => s(7)(131),lamdaOut => P(6)(267));
U_G7268: entity G port map(lamdaA => P(7)(260),lamdaB => P(7)(268),s => s(7)(132),lamdaOut => P(6)(268));
U_G7269: entity G port map(lamdaA => P(7)(261),lamdaB => P(7)(269),s => s(7)(133),lamdaOut => P(6)(269));
U_G7270: entity G port map(lamdaA => P(7)(262),lamdaB => P(7)(270),s => s(7)(134),lamdaOut => P(6)(270));
U_G7271: entity G port map(lamdaA => P(7)(263),lamdaB => P(7)(271),s => s(7)(135),lamdaOut => P(6)(271));
U_F7272: entity F port map(lamdaA => P(7)(272),lamdaB => P(7)(280),lamdaOut => P(6)(272));
U_F7273: entity F port map(lamdaA => P(7)(273),lamdaB => P(7)(281),lamdaOut => P(6)(273));
U_F7274: entity F port map(lamdaA => P(7)(274),lamdaB => P(7)(282),lamdaOut => P(6)(274));
U_F7275: entity F port map(lamdaA => P(7)(275),lamdaB => P(7)(283),lamdaOut => P(6)(275));
U_F7276: entity F port map(lamdaA => P(7)(276),lamdaB => P(7)(284),lamdaOut => P(6)(276));
U_F7277: entity F port map(lamdaA => P(7)(277),lamdaB => P(7)(285),lamdaOut => P(6)(277));
U_F7278: entity F port map(lamdaA => P(7)(278),lamdaB => P(7)(286),lamdaOut => P(6)(278));
U_F7279: entity F port map(lamdaA => P(7)(279),lamdaB => P(7)(287),lamdaOut => P(6)(279));
U_G7280: entity G port map(lamdaA => P(7)(272),lamdaB => P(7)(280),s => s(7)(136),lamdaOut => P(6)(280));
U_G7281: entity G port map(lamdaA => P(7)(273),lamdaB => P(7)(281),s => s(7)(137),lamdaOut => P(6)(281));
U_G7282: entity G port map(lamdaA => P(7)(274),lamdaB => P(7)(282),s => s(7)(138),lamdaOut => P(6)(282));
U_G7283: entity G port map(lamdaA => P(7)(275),lamdaB => P(7)(283),s => s(7)(139),lamdaOut => P(6)(283));
U_G7284: entity G port map(lamdaA => P(7)(276),lamdaB => P(7)(284),s => s(7)(140),lamdaOut => P(6)(284));
U_G7285: entity G port map(lamdaA => P(7)(277),lamdaB => P(7)(285),s => s(7)(141),lamdaOut => P(6)(285));
U_G7286: entity G port map(lamdaA => P(7)(278),lamdaB => P(7)(286),s => s(7)(142),lamdaOut => P(6)(286));
U_G7287: entity G port map(lamdaA => P(7)(279),lamdaB => P(7)(287),s => s(7)(143),lamdaOut => P(6)(287));
U_F7288: entity F port map(lamdaA => P(7)(288),lamdaB => P(7)(296),lamdaOut => P(6)(288));
U_F7289: entity F port map(lamdaA => P(7)(289),lamdaB => P(7)(297),lamdaOut => P(6)(289));
U_F7290: entity F port map(lamdaA => P(7)(290),lamdaB => P(7)(298),lamdaOut => P(6)(290));
U_F7291: entity F port map(lamdaA => P(7)(291),lamdaB => P(7)(299),lamdaOut => P(6)(291));
U_F7292: entity F port map(lamdaA => P(7)(292),lamdaB => P(7)(300),lamdaOut => P(6)(292));
U_F7293: entity F port map(lamdaA => P(7)(293),lamdaB => P(7)(301),lamdaOut => P(6)(293));
U_F7294: entity F port map(lamdaA => P(7)(294),lamdaB => P(7)(302),lamdaOut => P(6)(294));
U_F7295: entity F port map(lamdaA => P(7)(295),lamdaB => P(7)(303),lamdaOut => P(6)(295));
U_G7296: entity G port map(lamdaA => P(7)(288),lamdaB => P(7)(296),s => s(7)(144),lamdaOut => P(6)(296));
U_G7297: entity G port map(lamdaA => P(7)(289),lamdaB => P(7)(297),s => s(7)(145),lamdaOut => P(6)(297));
U_G7298: entity G port map(lamdaA => P(7)(290),lamdaB => P(7)(298),s => s(7)(146),lamdaOut => P(6)(298));
U_G7299: entity G port map(lamdaA => P(7)(291),lamdaB => P(7)(299),s => s(7)(147),lamdaOut => P(6)(299));
U_G7300: entity G port map(lamdaA => P(7)(292),lamdaB => P(7)(300),s => s(7)(148),lamdaOut => P(6)(300));
U_G7301: entity G port map(lamdaA => P(7)(293),lamdaB => P(7)(301),s => s(7)(149),lamdaOut => P(6)(301));
U_G7302: entity G port map(lamdaA => P(7)(294),lamdaB => P(7)(302),s => s(7)(150),lamdaOut => P(6)(302));
U_G7303: entity G port map(lamdaA => P(7)(295),lamdaB => P(7)(303),s => s(7)(151),lamdaOut => P(6)(303));
U_F7304: entity F port map(lamdaA => P(7)(304),lamdaB => P(7)(312),lamdaOut => P(6)(304));
U_F7305: entity F port map(lamdaA => P(7)(305),lamdaB => P(7)(313),lamdaOut => P(6)(305));
U_F7306: entity F port map(lamdaA => P(7)(306),lamdaB => P(7)(314),lamdaOut => P(6)(306));
U_F7307: entity F port map(lamdaA => P(7)(307),lamdaB => P(7)(315),lamdaOut => P(6)(307));
U_F7308: entity F port map(lamdaA => P(7)(308),lamdaB => P(7)(316),lamdaOut => P(6)(308));
U_F7309: entity F port map(lamdaA => P(7)(309),lamdaB => P(7)(317),lamdaOut => P(6)(309));
U_F7310: entity F port map(lamdaA => P(7)(310),lamdaB => P(7)(318),lamdaOut => P(6)(310));
U_F7311: entity F port map(lamdaA => P(7)(311),lamdaB => P(7)(319),lamdaOut => P(6)(311));
U_G7312: entity G port map(lamdaA => P(7)(304),lamdaB => P(7)(312),s => s(7)(152),lamdaOut => P(6)(312));
U_G7313: entity G port map(lamdaA => P(7)(305),lamdaB => P(7)(313),s => s(7)(153),lamdaOut => P(6)(313));
U_G7314: entity G port map(lamdaA => P(7)(306),lamdaB => P(7)(314),s => s(7)(154),lamdaOut => P(6)(314));
U_G7315: entity G port map(lamdaA => P(7)(307),lamdaB => P(7)(315),s => s(7)(155),lamdaOut => P(6)(315));
U_G7316: entity G port map(lamdaA => P(7)(308),lamdaB => P(7)(316),s => s(7)(156),lamdaOut => P(6)(316));
U_G7317: entity G port map(lamdaA => P(7)(309),lamdaB => P(7)(317),s => s(7)(157),lamdaOut => P(6)(317));
U_G7318: entity G port map(lamdaA => P(7)(310),lamdaB => P(7)(318),s => s(7)(158),lamdaOut => P(6)(318));
U_G7319: entity G port map(lamdaA => P(7)(311),lamdaB => P(7)(319),s => s(7)(159),lamdaOut => P(6)(319));
U_F7320: entity F port map(lamdaA => P(7)(320),lamdaB => P(7)(328),lamdaOut => P(6)(320));
U_F7321: entity F port map(lamdaA => P(7)(321),lamdaB => P(7)(329),lamdaOut => P(6)(321));
U_F7322: entity F port map(lamdaA => P(7)(322),lamdaB => P(7)(330),lamdaOut => P(6)(322));
U_F7323: entity F port map(lamdaA => P(7)(323),lamdaB => P(7)(331),lamdaOut => P(6)(323));
U_F7324: entity F port map(lamdaA => P(7)(324),lamdaB => P(7)(332),lamdaOut => P(6)(324));
U_F7325: entity F port map(lamdaA => P(7)(325),lamdaB => P(7)(333),lamdaOut => P(6)(325));
U_F7326: entity F port map(lamdaA => P(7)(326),lamdaB => P(7)(334),lamdaOut => P(6)(326));
U_F7327: entity F port map(lamdaA => P(7)(327),lamdaB => P(7)(335),lamdaOut => P(6)(327));
U_G7328: entity G port map(lamdaA => P(7)(320),lamdaB => P(7)(328),s => s(7)(160),lamdaOut => P(6)(328));
U_G7329: entity G port map(lamdaA => P(7)(321),lamdaB => P(7)(329),s => s(7)(161),lamdaOut => P(6)(329));
U_G7330: entity G port map(lamdaA => P(7)(322),lamdaB => P(7)(330),s => s(7)(162),lamdaOut => P(6)(330));
U_G7331: entity G port map(lamdaA => P(7)(323),lamdaB => P(7)(331),s => s(7)(163),lamdaOut => P(6)(331));
U_G7332: entity G port map(lamdaA => P(7)(324),lamdaB => P(7)(332),s => s(7)(164),lamdaOut => P(6)(332));
U_G7333: entity G port map(lamdaA => P(7)(325),lamdaB => P(7)(333),s => s(7)(165),lamdaOut => P(6)(333));
U_G7334: entity G port map(lamdaA => P(7)(326),lamdaB => P(7)(334),s => s(7)(166),lamdaOut => P(6)(334));
U_G7335: entity G port map(lamdaA => P(7)(327),lamdaB => P(7)(335),s => s(7)(167),lamdaOut => P(6)(335));
U_F7336: entity F port map(lamdaA => P(7)(336),lamdaB => P(7)(344),lamdaOut => P(6)(336));
U_F7337: entity F port map(lamdaA => P(7)(337),lamdaB => P(7)(345),lamdaOut => P(6)(337));
U_F7338: entity F port map(lamdaA => P(7)(338),lamdaB => P(7)(346),lamdaOut => P(6)(338));
U_F7339: entity F port map(lamdaA => P(7)(339),lamdaB => P(7)(347),lamdaOut => P(6)(339));
U_F7340: entity F port map(lamdaA => P(7)(340),lamdaB => P(7)(348),lamdaOut => P(6)(340));
U_F7341: entity F port map(lamdaA => P(7)(341),lamdaB => P(7)(349),lamdaOut => P(6)(341));
U_F7342: entity F port map(lamdaA => P(7)(342),lamdaB => P(7)(350),lamdaOut => P(6)(342));
U_F7343: entity F port map(lamdaA => P(7)(343),lamdaB => P(7)(351),lamdaOut => P(6)(343));
U_G7344: entity G port map(lamdaA => P(7)(336),lamdaB => P(7)(344),s => s(7)(168),lamdaOut => P(6)(344));
U_G7345: entity G port map(lamdaA => P(7)(337),lamdaB => P(7)(345),s => s(7)(169),lamdaOut => P(6)(345));
U_G7346: entity G port map(lamdaA => P(7)(338),lamdaB => P(7)(346),s => s(7)(170),lamdaOut => P(6)(346));
U_G7347: entity G port map(lamdaA => P(7)(339),lamdaB => P(7)(347),s => s(7)(171),lamdaOut => P(6)(347));
U_G7348: entity G port map(lamdaA => P(7)(340),lamdaB => P(7)(348),s => s(7)(172),lamdaOut => P(6)(348));
U_G7349: entity G port map(lamdaA => P(7)(341),lamdaB => P(7)(349),s => s(7)(173),lamdaOut => P(6)(349));
U_G7350: entity G port map(lamdaA => P(7)(342),lamdaB => P(7)(350),s => s(7)(174),lamdaOut => P(6)(350));
U_G7351: entity G port map(lamdaA => P(7)(343),lamdaB => P(7)(351),s => s(7)(175),lamdaOut => P(6)(351));
U_F7352: entity F port map(lamdaA => P(7)(352),lamdaB => P(7)(360),lamdaOut => P(6)(352));
U_F7353: entity F port map(lamdaA => P(7)(353),lamdaB => P(7)(361),lamdaOut => P(6)(353));
U_F7354: entity F port map(lamdaA => P(7)(354),lamdaB => P(7)(362),lamdaOut => P(6)(354));
U_F7355: entity F port map(lamdaA => P(7)(355),lamdaB => P(7)(363),lamdaOut => P(6)(355));
U_F7356: entity F port map(lamdaA => P(7)(356),lamdaB => P(7)(364),lamdaOut => P(6)(356));
U_F7357: entity F port map(lamdaA => P(7)(357),lamdaB => P(7)(365),lamdaOut => P(6)(357));
U_F7358: entity F port map(lamdaA => P(7)(358),lamdaB => P(7)(366),lamdaOut => P(6)(358));
U_F7359: entity F port map(lamdaA => P(7)(359),lamdaB => P(7)(367),lamdaOut => P(6)(359));
U_G7360: entity G port map(lamdaA => P(7)(352),lamdaB => P(7)(360),s => s(7)(176),lamdaOut => P(6)(360));
U_G7361: entity G port map(lamdaA => P(7)(353),lamdaB => P(7)(361),s => s(7)(177),lamdaOut => P(6)(361));
U_G7362: entity G port map(lamdaA => P(7)(354),lamdaB => P(7)(362),s => s(7)(178),lamdaOut => P(6)(362));
U_G7363: entity G port map(lamdaA => P(7)(355),lamdaB => P(7)(363),s => s(7)(179),lamdaOut => P(6)(363));
U_G7364: entity G port map(lamdaA => P(7)(356),lamdaB => P(7)(364),s => s(7)(180),lamdaOut => P(6)(364));
U_G7365: entity G port map(lamdaA => P(7)(357),lamdaB => P(7)(365),s => s(7)(181),lamdaOut => P(6)(365));
U_G7366: entity G port map(lamdaA => P(7)(358),lamdaB => P(7)(366),s => s(7)(182),lamdaOut => P(6)(366));
U_G7367: entity G port map(lamdaA => P(7)(359),lamdaB => P(7)(367),s => s(7)(183),lamdaOut => P(6)(367));
U_F7368: entity F port map(lamdaA => P(7)(368),lamdaB => P(7)(376),lamdaOut => P(6)(368));
U_F7369: entity F port map(lamdaA => P(7)(369),lamdaB => P(7)(377),lamdaOut => P(6)(369));
U_F7370: entity F port map(lamdaA => P(7)(370),lamdaB => P(7)(378),lamdaOut => P(6)(370));
U_F7371: entity F port map(lamdaA => P(7)(371),lamdaB => P(7)(379),lamdaOut => P(6)(371));
U_F7372: entity F port map(lamdaA => P(7)(372),lamdaB => P(7)(380),lamdaOut => P(6)(372));
U_F7373: entity F port map(lamdaA => P(7)(373),lamdaB => P(7)(381),lamdaOut => P(6)(373));
U_F7374: entity F port map(lamdaA => P(7)(374),lamdaB => P(7)(382),lamdaOut => P(6)(374));
U_F7375: entity F port map(lamdaA => P(7)(375),lamdaB => P(7)(383),lamdaOut => P(6)(375));
U_G7376: entity G port map(lamdaA => P(7)(368),lamdaB => P(7)(376),s => s(7)(184),lamdaOut => P(6)(376));
U_G7377: entity G port map(lamdaA => P(7)(369),lamdaB => P(7)(377),s => s(7)(185),lamdaOut => P(6)(377));
U_G7378: entity G port map(lamdaA => P(7)(370),lamdaB => P(7)(378),s => s(7)(186),lamdaOut => P(6)(378));
U_G7379: entity G port map(lamdaA => P(7)(371),lamdaB => P(7)(379),s => s(7)(187),lamdaOut => P(6)(379));
U_G7380: entity G port map(lamdaA => P(7)(372),lamdaB => P(7)(380),s => s(7)(188),lamdaOut => P(6)(380));
U_G7381: entity G port map(lamdaA => P(7)(373),lamdaB => P(7)(381),s => s(7)(189),lamdaOut => P(6)(381));
U_G7382: entity G port map(lamdaA => P(7)(374),lamdaB => P(7)(382),s => s(7)(190),lamdaOut => P(6)(382));
U_G7383: entity G port map(lamdaA => P(7)(375),lamdaB => P(7)(383),s => s(7)(191),lamdaOut => P(6)(383));
U_F7384: entity F port map(lamdaA => P(7)(384),lamdaB => P(7)(392),lamdaOut => P(6)(384));
U_F7385: entity F port map(lamdaA => P(7)(385),lamdaB => P(7)(393),lamdaOut => P(6)(385));
U_F7386: entity F port map(lamdaA => P(7)(386),lamdaB => P(7)(394),lamdaOut => P(6)(386));
U_F7387: entity F port map(lamdaA => P(7)(387),lamdaB => P(7)(395),lamdaOut => P(6)(387));
U_F7388: entity F port map(lamdaA => P(7)(388),lamdaB => P(7)(396),lamdaOut => P(6)(388));
U_F7389: entity F port map(lamdaA => P(7)(389),lamdaB => P(7)(397),lamdaOut => P(6)(389));
U_F7390: entity F port map(lamdaA => P(7)(390),lamdaB => P(7)(398),lamdaOut => P(6)(390));
U_F7391: entity F port map(lamdaA => P(7)(391),lamdaB => P(7)(399),lamdaOut => P(6)(391));
U_G7392: entity G port map(lamdaA => P(7)(384),lamdaB => P(7)(392),s => s(7)(192),lamdaOut => P(6)(392));
U_G7393: entity G port map(lamdaA => P(7)(385),lamdaB => P(7)(393),s => s(7)(193),lamdaOut => P(6)(393));
U_G7394: entity G port map(lamdaA => P(7)(386),lamdaB => P(7)(394),s => s(7)(194),lamdaOut => P(6)(394));
U_G7395: entity G port map(lamdaA => P(7)(387),lamdaB => P(7)(395),s => s(7)(195),lamdaOut => P(6)(395));
U_G7396: entity G port map(lamdaA => P(7)(388),lamdaB => P(7)(396),s => s(7)(196),lamdaOut => P(6)(396));
U_G7397: entity G port map(lamdaA => P(7)(389),lamdaB => P(7)(397),s => s(7)(197),lamdaOut => P(6)(397));
U_G7398: entity G port map(lamdaA => P(7)(390),lamdaB => P(7)(398),s => s(7)(198),lamdaOut => P(6)(398));
U_G7399: entity G port map(lamdaA => P(7)(391),lamdaB => P(7)(399),s => s(7)(199),lamdaOut => P(6)(399));
U_F7400: entity F port map(lamdaA => P(7)(400),lamdaB => P(7)(408),lamdaOut => P(6)(400));
U_F7401: entity F port map(lamdaA => P(7)(401),lamdaB => P(7)(409),lamdaOut => P(6)(401));
U_F7402: entity F port map(lamdaA => P(7)(402),lamdaB => P(7)(410),lamdaOut => P(6)(402));
U_F7403: entity F port map(lamdaA => P(7)(403),lamdaB => P(7)(411),lamdaOut => P(6)(403));
U_F7404: entity F port map(lamdaA => P(7)(404),lamdaB => P(7)(412),lamdaOut => P(6)(404));
U_F7405: entity F port map(lamdaA => P(7)(405),lamdaB => P(7)(413),lamdaOut => P(6)(405));
U_F7406: entity F port map(lamdaA => P(7)(406),lamdaB => P(7)(414),lamdaOut => P(6)(406));
U_F7407: entity F port map(lamdaA => P(7)(407),lamdaB => P(7)(415),lamdaOut => P(6)(407));
U_G7408: entity G port map(lamdaA => P(7)(400),lamdaB => P(7)(408),s => s(7)(200),lamdaOut => P(6)(408));
U_G7409: entity G port map(lamdaA => P(7)(401),lamdaB => P(7)(409),s => s(7)(201),lamdaOut => P(6)(409));
U_G7410: entity G port map(lamdaA => P(7)(402),lamdaB => P(7)(410),s => s(7)(202),lamdaOut => P(6)(410));
U_G7411: entity G port map(lamdaA => P(7)(403),lamdaB => P(7)(411),s => s(7)(203),lamdaOut => P(6)(411));
U_G7412: entity G port map(lamdaA => P(7)(404),lamdaB => P(7)(412),s => s(7)(204),lamdaOut => P(6)(412));
U_G7413: entity G port map(lamdaA => P(7)(405),lamdaB => P(7)(413),s => s(7)(205),lamdaOut => P(6)(413));
U_G7414: entity G port map(lamdaA => P(7)(406),lamdaB => P(7)(414),s => s(7)(206),lamdaOut => P(6)(414));
U_G7415: entity G port map(lamdaA => P(7)(407),lamdaB => P(7)(415),s => s(7)(207),lamdaOut => P(6)(415));
U_F7416: entity F port map(lamdaA => P(7)(416),lamdaB => P(7)(424),lamdaOut => P(6)(416));
U_F7417: entity F port map(lamdaA => P(7)(417),lamdaB => P(7)(425),lamdaOut => P(6)(417));
U_F7418: entity F port map(lamdaA => P(7)(418),lamdaB => P(7)(426),lamdaOut => P(6)(418));
U_F7419: entity F port map(lamdaA => P(7)(419),lamdaB => P(7)(427),lamdaOut => P(6)(419));
U_F7420: entity F port map(lamdaA => P(7)(420),lamdaB => P(7)(428),lamdaOut => P(6)(420));
U_F7421: entity F port map(lamdaA => P(7)(421),lamdaB => P(7)(429),lamdaOut => P(6)(421));
U_F7422: entity F port map(lamdaA => P(7)(422),lamdaB => P(7)(430),lamdaOut => P(6)(422));
U_F7423: entity F port map(lamdaA => P(7)(423),lamdaB => P(7)(431),lamdaOut => P(6)(423));
U_G7424: entity G port map(lamdaA => P(7)(416),lamdaB => P(7)(424),s => s(7)(208),lamdaOut => P(6)(424));
U_G7425: entity G port map(lamdaA => P(7)(417),lamdaB => P(7)(425),s => s(7)(209),lamdaOut => P(6)(425));
U_G7426: entity G port map(lamdaA => P(7)(418),lamdaB => P(7)(426),s => s(7)(210),lamdaOut => P(6)(426));
U_G7427: entity G port map(lamdaA => P(7)(419),lamdaB => P(7)(427),s => s(7)(211),lamdaOut => P(6)(427));
U_G7428: entity G port map(lamdaA => P(7)(420),lamdaB => P(7)(428),s => s(7)(212),lamdaOut => P(6)(428));
U_G7429: entity G port map(lamdaA => P(7)(421),lamdaB => P(7)(429),s => s(7)(213),lamdaOut => P(6)(429));
U_G7430: entity G port map(lamdaA => P(7)(422),lamdaB => P(7)(430),s => s(7)(214),lamdaOut => P(6)(430));
U_G7431: entity G port map(lamdaA => P(7)(423),lamdaB => P(7)(431),s => s(7)(215),lamdaOut => P(6)(431));
U_F7432: entity F port map(lamdaA => P(7)(432),lamdaB => P(7)(440),lamdaOut => P(6)(432));
U_F7433: entity F port map(lamdaA => P(7)(433),lamdaB => P(7)(441),lamdaOut => P(6)(433));
U_F7434: entity F port map(lamdaA => P(7)(434),lamdaB => P(7)(442),lamdaOut => P(6)(434));
U_F7435: entity F port map(lamdaA => P(7)(435),lamdaB => P(7)(443),lamdaOut => P(6)(435));
U_F7436: entity F port map(lamdaA => P(7)(436),lamdaB => P(7)(444),lamdaOut => P(6)(436));
U_F7437: entity F port map(lamdaA => P(7)(437),lamdaB => P(7)(445),lamdaOut => P(6)(437));
U_F7438: entity F port map(lamdaA => P(7)(438),lamdaB => P(7)(446),lamdaOut => P(6)(438));
U_F7439: entity F port map(lamdaA => P(7)(439),lamdaB => P(7)(447),lamdaOut => P(6)(439));
U_G7440: entity G port map(lamdaA => P(7)(432),lamdaB => P(7)(440),s => s(7)(216),lamdaOut => P(6)(440));
U_G7441: entity G port map(lamdaA => P(7)(433),lamdaB => P(7)(441),s => s(7)(217),lamdaOut => P(6)(441));
U_G7442: entity G port map(lamdaA => P(7)(434),lamdaB => P(7)(442),s => s(7)(218),lamdaOut => P(6)(442));
U_G7443: entity G port map(lamdaA => P(7)(435),lamdaB => P(7)(443),s => s(7)(219),lamdaOut => P(6)(443));
U_G7444: entity G port map(lamdaA => P(7)(436),lamdaB => P(7)(444),s => s(7)(220),lamdaOut => P(6)(444));
U_G7445: entity G port map(lamdaA => P(7)(437),lamdaB => P(7)(445),s => s(7)(221),lamdaOut => P(6)(445));
U_G7446: entity G port map(lamdaA => P(7)(438),lamdaB => P(7)(446),s => s(7)(222),lamdaOut => P(6)(446));
U_G7447: entity G port map(lamdaA => P(7)(439),lamdaB => P(7)(447),s => s(7)(223),lamdaOut => P(6)(447));
U_F7448: entity F port map(lamdaA => P(7)(448),lamdaB => P(7)(456),lamdaOut => P(6)(448));
U_F7449: entity F port map(lamdaA => P(7)(449),lamdaB => P(7)(457),lamdaOut => P(6)(449));
U_F7450: entity F port map(lamdaA => P(7)(450),lamdaB => P(7)(458),lamdaOut => P(6)(450));
U_F7451: entity F port map(lamdaA => P(7)(451),lamdaB => P(7)(459),lamdaOut => P(6)(451));
U_F7452: entity F port map(lamdaA => P(7)(452),lamdaB => P(7)(460),lamdaOut => P(6)(452));
U_F7453: entity F port map(lamdaA => P(7)(453),lamdaB => P(7)(461),lamdaOut => P(6)(453));
U_F7454: entity F port map(lamdaA => P(7)(454),lamdaB => P(7)(462),lamdaOut => P(6)(454));
U_F7455: entity F port map(lamdaA => P(7)(455),lamdaB => P(7)(463),lamdaOut => P(6)(455));
U_G7456: entity G port map(lamdaA => P(7)(448),lamdaB => P(7)(456),s => s(7)(224),lamdaOut => P(6)(456));
U_G7457: entity G port map(lamdaA => P(7)(449),lamdaB => P(7)(457),s => s(7)(225),lamdaOut => P(6)(457));
U_G7458: entity G port map(lamdaA => P(7)(450),lamdaB => P(7)(458),s => s(7)(226),lamdaOut => P(6)(458));
U_G7459: entity G port map(lamdaA => P(7)(451),lamdaB => P(7)(459),s => s(7)(227),lamdaOut => P(6)(459));
U_G7460: entity G port map(lamdaA => P(7)(452),lamdaB => P(7)(460),s => s(7)(228),lamdaOut => P(6)(460));
U_G7461: entity G port map(lamdaA => P(7)(453),lamdaB => P(7)(461),s => s(7)(229),lamdaOut => P(6)(461));
U_G7462: entity G port map(lamdaA => P(7)(454),lamdaB => P(7)(462),s => s(7)(230),lamdaOut => P(6)(462));
U_G7463: entity G port map(lamdaA => P(7)(455),lamdaB => P(7)(463),s => s(7)(231),lamdaOut => P(6)(463));
U_F7464: entity F port map(lamdaA => P(7)(464),lamdaB => P(7)(472),lamdaOut => P(6)(464));
U_F7465: entity F port map(lamdaA => P(7)(465),lamdaB => P(7)(473),lamdaOut => P(6)(465));
U_F7466: entity F port map(lamdaA => P(7)(466),lamdaB => P(7)(474),lamdaOut => P(6)(466));
U_F7467: entity F port map(lamdaA => P(7)(467),lamdaB => P(7)(475),lamdaOut => P(6)(467));
U_F7468: entity F port map(lamdaA => P(7)(468),lamdaB => P(7)(476),lamdaOut => P(6)(468));
U_F7469: entity F port map(lamdaA => P(7)(469),lamdaB => P(7)(477),lamdaOut => P(6)(469));
U_F7470: entity F port map(lamdaA => P(7)(470),lamdaB => P(7)(478),lamdaOut => P(6)(470));
U_F7471: entity F port map(lamdaA => P(7)(471),lamdaB => P(7)(479),lamdaOut => P(6)(471));
U_G7472: entity G port map(lamdaA => P(7)(464),lamdaB => P(7)(472),s => s(7)(232),lamdaOut => P(6)(472));
U_G7473: entity G port map(lamdaA => P(7)(465),lamdaB => P(7)(473),s => s(7)(233),lamdaOut => P(6)(473));
U_G7474: entity G port map(lamdaA => P(7)(466),lamdaB => P(7)(474),s => s(7)(234),lamdaOut => P(6)(474));
U_G7475: entity G port map(lamdaA => P(7)(467),lamdaB => P(7)(475),s => s(7)(235),lamdaOut => P(6)(475));
U_G7476: entity G port map(lamdaA => P(7)(468),lamdaB => P(7)(476),s => s(7)(236),lamdaOut => P(6)(476));
U_G7477: entity G port map(lamdaA => P(7)(469),lamdaB => P(7)(477),s => s(7)(237),lamdaOut => P(6)(477));
U_G7478: entity G port map(lamdaA => P(7)(470),lamdaB => P(7)(478),s => s(7)(238),lamdaOut => P(6)(478));
U_G7479: entity G port map(lamdaA => P(7)(471),lamdaB => P(7)(479),s => s(7)(239),lamdaOut => P(6)(479));
U_F7480: entity F port map(lamdaA => P(7)(480),lamdaB => P(7)(488),lamdaOut => P(6)(480));
U_F7481: entity F port map(lamdaA => P(7)(481),lamdaB => P(7)(489),lamdaOut => P(6)(481));
U_F7482: entity F port map(lamdaA => P(7)(482),lamdaB => P(7)(490),lamdaOut => P(6)(482));
U_F7483: entity F port map(lamdaA => P(7)(483),lamdaB => P(7)(491),lamdaOut => P(6)(483));
U_F7484: entity F port map(lamdaA => P(7)(484),lamdaB => P(7)(492),lamdaOut => P(6)(484));
U_F7485: entity F port map(lamdaA => P(7)(485),lamdaB => P(7)(493),lamdaOut => P(6)(485));
U_F7486: entity F port map(lamdaA => P(7)(486),lamdaB => P(7)(494),lamdaOut => P(6)(486));
U_F7487: entity F port map(lamdaA => P(7)(487),lamdaB => P(7)(495),lamdaOut => P(6)(487));
U_G7488: entity G port map(lamdaA => P(7)(480),lamdaB => P(7)(488),s => s(7)(240),lamdaOut => P(6)(488));
U_G7489: entity G port map(lamdaA => P(7)(481),lamdaB => P(7)(489),s => s(7)(241),lamdaOut => P(6)(489));
U_G7490: entity G port map(lamdaA => P(7)(482),lamdaB => P(7)(490),s => s(7)(242),lamdaOut => P(6)(490));
U_G7491: entity G port map(lamdaA => P(7)(483),lamdaB => P(7)(491),s => s(7)(243),lamdaOut => P(6)(491));
U_G7492: entity G port map(lamdaA => P(7)(484),lamdaB => P(7)(492),s => s(7)(244),lamdaOut => P(6)(492));
U_G7493: entity G port map(lamdaA => P(7)(485),lamdaB => P(7)(493),s => s(7)(245),lamdaOut => P(6)(493));
U_G7494: entity G port map(lamdaA => P(7)(486),lamdaB => P(7)(494),s => s(7)(246),lamdaOut => P(6)(494));
U_G7495: entity G port map(lamdaA => P(7)(487),lamdaB => P(7)(495),s => s(7)(247),lamdaOut => P(6)(495));
U_F7496: entity F port map(lamdaA => P(7)(496),lamdaB => P(7)(504),lamdaOut => P(6)(496));
U_F7497: entity F port map(lamdaA => P(7)(497),lamdaB => P(7)(505),lamdaOut => P(6)(497));
U_F7498: entity F port map(lamdaA => P(7)(498),lamdaB => P(7)(506),lamdaOut => P(6)(498));
U_F7499: entity F port map(lamdaA => P(7)(499),lamdaB => P(7)(507),lamdaOut => P(6)(499));
U_F7500: entity F port map(lamdaA => P(7)(500),lamdaB => P(7)(508),lamdaOut => P(6)(500));
U_F7501: entity F port map(lamdaA => P(7)(501),lamdaB => P(7)(509),lamdaOut => P(6)(501));
U_F7502: entity F port map(lamdaA => P(7)(502),lamdaB => P(7)(510),lamdaOut => P(6)(502));
U_F7503: entity F port map(lamdaA => P(7)(503),lamdaB => P(7)(511),lamdaOut => P(6)(503));
U_G7504: entity G port map(lamdaA => P(7)(496),lamdaB => P(7)(504),s => s(7)(248),lamdaOut => P(6)(504));
U_G7505: entity G port map(lamdaA => P(7)(497),lamdaB => P(7)(505),s => s(7)(249),lamdaOut => P(6)(505));
U_G7506: entity G port map(lamdaA => P(7)(498),lamdaB => P(7)(506),s => s(7)(250),lamdaOut => P(6)(506));
U_G7507: entity G port map(lamdaA => P(7)(499),lamdaB => P(7)(507),s => s(7)(251),lamdaOut => P(6)(507));
U_G7508: entity G port map(lamdaA => P(7)(500),lamdaB => P(7)(508),s => s(7)(252),lamdaOut => P(6)(508));
U_G7509: entity G port map(lamdaA => P(7)(501),lamdaB => P(7)(509),s => s(7)(253),lamdaOut => P(6)(509));
U_G7510: entity G port map(lamdaA => P(7)(502),lamdaB => P(7)(510),s => s(7)(254),lamdaOut => P(6)(510));
U_G7511: entity G port map(lamdaA => P(7)(503),lamdaB => P(7)(511),s => s(7)(255),lamdaOut => P(6)(511));
U_F7512: entity F port map(lamdaA => P(7)(512),lamdaB => P(7)(520),lamdaOut => P(6)(512));
U_F7513: entity F port map(lamdaA => P(7)(513),lamdaB => P(7)(521),lamdaOut => P(6)(513));
U_F7514: entity F port map(lamdaA => P(7)(514),lamdaB => P(7)(522),lamdaOut => P(6)(514));
U_F7515: entity F port map(lamdaA => P(7)(515),lamdaB => P(7)(523),lamdaOut => P(6)(515));
U_F7516: entity F port map(lamdaA => P(7)(516),lamdaB => P(7)(524),lamdaOut => P(6)(516));
U_F7517: entity F port map(lamdaA => P(7)(517),lamdaB => P(7)(525),lamdaOut => P(6)(517));
U_F7518: entity F port map(lamdaA => P(7)(518),lamdaB => P(7)(526),lamdaOut => P(6)(518));
U_F7519: entity F port map(lamdaA => P(7)(519),lamdaB => P(7)(527),lamdaOut => P(6)(519));
U_G7520: entity G port map(lamdaA => P(7)(512),lamdaB => P(7)(520),s => s(7)(256),lamdaOut => P(6)(520));
U_G7521: entity G port map(lamdaA => P(7)(513),lamdaB => P(7)(521),s => s(7)(257),lamdaOut => P(6)(521));
U_G7522: entity G port map(lamdaA => P(7)(514),lamdaB => P(7)(522),s => s(7)(258),lamdaOut => P(6)(522));
U_G7523: entity G port map(lamdaA => P(7)(515),lamdaB => P(7)(523),s => s(7)(259),lamdaOut => P(6)(523));
U_G7524: entity G port map(lamdaA => P(7)(516),lamdaB => P(7)(524),s => s(7)(260),lamdaOut => P(6)(524));
U_G7525: entity G port map(lamdaA => P(7)(517),lamdaB => P(7)(525),s => s(7)(261),lamdaOut => P(6)(525));
U_G7526: entity G port map(lamdaA => P(7)(518),lamdaB => P(7)(526),s => s(7)(262),lamdaOut => P(6)(526));
U_G7527: entity G port map(lamdaA => P(7)(519),lamdaB => P(7)(527),s => s(7)(263),lamdaOut => P(6)(527));
U_F7528: entity F port map(lamdaA => P(7)(528),lamdaB => P(7)(536),lamdaOut => P(6)(528));
U_F7529: entity F port map(lamdaA => P(7)(529),lamdaB => P(7)(537),lamdaOut => P(6)(529));
U_F7530: entity F port map(lamdaA => P(7)(530),lamdaB => P(7)(538),lamdaOut => P(6)(530));
U_F7531: entity F port map(lamdaA => P(7)(531),lamdaB => P(7)(539),lamdaOut => P(6)(531));
U_F7532: entity F port map(lamdaA => P(7)(532),lamdaB => P(7)(540),lamdaOut => P(6)(532));
U_F7533: entity F port map(lamdaA => P(7)(533),lamdaB => P(7)(541),lamdaOut => P(6)(533));
U_F7534: entity F port map(lamdaA => P(7)(534),lamdaB => P(7)(542),lamdaOut => P(6)(534));
U_F7535: entity F port map(lamdaA => P(7)(535),lamdaB => P(7)(543),lamdaOut => P(6)(535));
U_G7536: entity G port map(lamdaA => P(7)(528),lamdaB => P(7)(536),s => s(7)(264),lamdaOut => P(6)(536));
U_G7537: entity G port map(lamdaA => P(7)(529),lamdaB => P(7)(537),s => s(7)(265),lamdaOut => P(6)(537));
U_G7538: entity G port map(lamdaA => P(7)(530),lamdaB => P(7)(538),s => s(7)(266),lamdaOut => P(6)(538));
U_G7539: entity G port map(lamdaA => P(7)(531),lamdaB => P(7)(539),s => s(7)(267),lamdaOut => P(6)(539));
U_G7540: entity G port map(lamdaA => P(7)(532),lamdaB => P(7)(540),s => s(7)(268),lamdaOut => P(6)(540));
U_G7541: entity G port map(lamdaA => P(7)(533),lamdaB => P(7)(541),s => s(7)(269),lamdaOut => P(6)(541));
U_G7542: entity G port map(lamdaA => P(7)(534),lamdaB => P(7)(542),s => s(7)(270),lamdaOut => P(6)(542));
U_G7543: entity G port map(lamdaA => P(7)(535),lamdaB => P(7)(543),s => s(7)(271),lamdaOut => P(6)(543));
U_F7544: entity F port map(lamdaA => P(7)(544),lamdaB => P(7)(552),lamdaOut => P(6)(544));
U_F7545: entity F port map(lamdaA => P(7)(545),lamdaB => P(7)(553),lamdaOut => P(6)(545));
U_F7546: entity F port map(lamdaA => P(7)(546),lamdaB => P(7)(554),lamdaOut => P(6)(546));
U_F7547: entity F port map(lamdaA => P(7)(547),lamdaB => P(7)(555),lamdaOut => P(6)(547));
U_F7548: entity F port map(lamdaA => P(7)(548),lamdaB => P(7)(556),lamdaOut => P(6)(548));
U_F7549: entity F port map(lamdaA => P(7)(549),lamdaB => P(7)(557),lamdaOut => P(6)(549));
U_F7550: entity F port map(lamdaA => P(7)(550),lamdaB => P(7)(558),lamdaOut => P(6)(550));
U_F7551: entity F port map(lamdaA => P(7)(551),lamdaB => P(7)(559),lamdaOut => P(6)(551));
U_G7552: entity G port map(lamdaA => P(7)(544),lamdaB => P(7)(552),s => s(7)(272),lamdaOut => P(6)(552));
U_G7553: entity G port map(lamdaA => P(7)(545),lamdaB => P(7)(553),s => s(7)(273),lamdaOut => P(6)(553));
U_G7554: entity G port map(lamdaA => P(7)(546),lamdaB => P(7)(554),s => s(7)(274),lamdaOut => P(6)(554));
U_G7555: entity G port map(lamdaA => P(7)(547),lamdaB => P(7)(555),s => s(7)(275),lamdaOut => P(6)(555));
U_G7556: entity G port map(lamdaA => P(7)(548),lamdaB => P(7)(556),s => s(7)(276),lamdaOut => P(6)(556));
U_G7557: entity G port map(lamdaA => P(7)(549),lamdaB => P(7)(557),s => s(7)(277),lamdaOut => P(6)(557));
U_G7558: entity G port map(lamdaA => P(7)(550),lamdaB => P(7)(558),s => s(7)(278),lamdaOut => P(6)(558));
U_G7559: entity G port map(lamdaA => P(7)(551),lamdaB => P(7)(559),s => s(7)(279),lamdaOut => P(6)(559));
U_F7560: entity F port map(lamdaA => P(7)(560),lamdaB => P(7)(568),lamdaOut => P(6)(560));
U_F7561: entity F port map(lamdaA => P(7)(561),lamdaB => P(7)(569),lamdaOut => P(6)(561));
U_F7562: entity F port map(lamdaA => P(7)(562),lamdaB => P(7)(570),lamdaOut => P(6)(562));
U_F7563: entity F port map(lamdaA => P(7)(563),lamdaB => P(7)(571),lamdaOut => P(6)(563));
U_F7564: entity F port map(lamdaA => P(7)(564),lamdaB => P(7)(572),lamdaOut => P(6)(564));
U_F7565: entity F port map(lamdaA => P(7)(565),lamdaB => P(7)(573),lamdaOut => P(6)(565));
U_F7566: entity F port map(lamdaA => P(7)(566),lamdaB => P(7)(574),lamdaOut => P(6)(566));
U_F7567: entity F port map(lamdaA => P(7)(567),lamdaB => P(7)(575),lamdaOut => P(6)(567));
U_G7568: entity G port map(lamdaA => P(7)(560),lamdaB => P(7)(568),s => s(7)(280),lamdaOut => P(6)(568));
U_G7569: entity G port map(lamdaA => P(7)(561),lamdaB => P(7)(569),s => s(7)(281),lamdaOut => P(6)(569));
U_G7570: entity G port map(lamdaA => P(7)(562),lamdaB => P(7)(570),s => s(7)(282),lamdaOut => P(6)(570));
U_G7571: entity G port map(lamdaA => P(7)(563),lamdaB => P(7)(571),s => s(7)(283),lamdaOut => P(6)(571));
U_G7572: entity G port map(lamdaA => P(7)(564),lamdaB => P(7)(572),s => s(7)(284),lamdaOut => P(6)(572));
U_G7573: entity G port map(lamdaA => P(7)(565),lamdaB => P(7)(573),s => s(7)(285),lamdaOut => P(6)(573));
U_G7574: entity G port map(lamdaA => P(7)(566),lamdaB => P(7)(574),s => s(7)(286),lamdaOut => P(6)(574));
U_G7575: entity G port map(lamdaA => P(7)(567),lamdaB => P(7)(575),s => s(7)(287),lamdaOut => P(6)(575));
U_F7576: entity F port map(lamdaA => P(7)(576),lamdaB => P(7)(584),lamdaOut => P(6)(576));
U_F7577: entity F port map(lamdaA => P(7)(577),lamdaB => P(7)(585),lamdaOut => P(6)(577));
U_F7578: entity F port map(lamdaA => P(7)(578),lamdaB => P(7)(586),lamdaOut => P(6)(578));
U_F7579: entity F port map(lamdaA => P(7)(579),lamdaB => P(7)(587),lamdaOut => P(6)(579));
U_F7580: entity F port map(lamdaA => P(7)(580),lamdaB => P(7)(588),lamdaOut => P(6)(580));
U_F7581: entity F port map(lamdaA => P(7)(581),lamdaB => P(7)(589),lamdaOut => P(6)(581));
U_F7582: entity F port map(lamdaA => P(7)(582),lamdaB => P(7)(590),lamdaOut => P(6)(582));
U_F7583: entity F port map(lamdaA => P(7)(583),lamdaB => P(7)(591),lamdaOut => P(6)(583));
U_G7584: entity G port map(lamdaA => P(7)(576),lamdaB => P(7)(584),s => s(7)(288),lamdaOut => P(6)(584));
U_G7585: entity G port map(lamdaA => P(7)(577),lamdaB => P(7)(585),s => s(7)(289),lamdaOut => P(6)(585));
U_G7586: entity G port map(lamdaA => P(7)(578),lamdaB => P(7)(586),s => s(7)(290),lamdaOut => P(6)(586));
U_G7587: entity G port map(lamdaA => P(7)(579),lamdaB => P(7)(587),s => s(7)(291),lamdaOut => P(6)(587));
U_G7588: entity G port map(lamdaA => P(7)(580),lamdaB => P(7)(588),s => s(7)(292),lamdaOut => P(6)(588));
U_G7589: entity G port map(lamdaA => P(7)(581),lamdaB => P(7)(589),s => s(7)(293),lamdaOut => P(6)(589));
U_G7590: entity G port map(lamdaA => P(7)(582),lamdaB => P(7)(590),s => s(7)(294),lamdaOut => P(6)(590));
U_G7591: entity G port map(lamdaA => P(7)(583),lamdaB => P(7)(591),s => s(7)(295),lamdaOut => P(6)(591));
U_F7592: entity F port map(lamdaA => P(7)(592),lamdaB => P(7)(600),lamdaOut => P(6)(592));
U_F7593: entity F port map(lamdaA => P(7)(593),lamdaB => P(7)(601),lamdaOut => P(6)(593));
U_F7594: entity F port map(lamdaA => P(7)(594),lamdaB => P(7)(602),lamdaOut => P(6)(594));
U_F7595: entity F port map(lamdaA => P(7)(595),lamdaB => P(7)(603),lamdaOut => P(6)(595));
U_F7596: entity F port map(lamdaA => P(7)(596),lamdaB => P(7)(604),lamdaOut => P(6)(596));
U_F7597: entity F port map(lamdaA => P(7)(597),lamdaB => P(7)(605),lamdaOut => P(6)(597));
U_F7598: entity F port map(lamdaA => P(7)(598),lamdaB => P(7)(606),lamdaOut => P(6)(598));
U_F7599: entity F port map(lamdaA => P(7)(599),lamdaB => P(7)(607),lamdaOut => P(6)(599));
U_G7600: entity G port map(lamdaA => P(7)(592),lamdaB => P(7)(600),s => s(7)(296),lamdaOut => P(6)(600));
U_G7601: entity G port map(lamdaA => P(7)(593),lamdaB => P(7)(601),s => s(7)(297),lamdaOut => P(6)(601));
U_G7602: entity G port map(lamdaA => P(7)(594),lamdaB => P(7)(602),s => s(7)(298),lamdaOut => P(6)(602));
U_G7603: entity G port map(lamdaA => P(7)(595),lamdaB => P(7)(603),s => s(7)(299),lamdaOut => P(6)(603));
U_G7604: entity G port map(lamdaA => P(7)(596),lamdaB => P(7)(604),s => s(7)(300),lamdaOut => P(6)(604));
U_G7605: entity G port map(lamdaA => P(7)(597),lamdaB => P(7)(605),s => s(7)(301),lamdaOut => P(6)(605));
U_G7606: entity G port map(lamdaA => P(7)(598),lamdaB => P(7)(606),s => s(7)(302),lamdaOut => P(6)(606));
U_G7607: entity G port map(lamdaA => P(7)(599),lamdaB => P(7)(607),s => s(7)(303),lamdaOut => P(6)(607));
U_F7608: entity F port map(lamdaA => P(7)(608),lamdaB => P(7)(616),lamdaOut => P(6)(608));
U_F7609: entity F port map(lamdaA => P(7)(609),lamdaB => P(7)(617),lamdaOut => P(6)(609));
U_F7610: entity F port map(lamdaA => P(7)(610),lamdaB => P(7)(618),lamdaOut => P(6)(610));
U_F7611: entity F port map(lamdaA => P(7)(611),lamdaB => P(7)(619),lamdaOut => P(6)(611));
U_F7612: entity F port map(lamdaA => P(7)(612),lamdaB => P(7)(620),lamdaOut => P(6)(612));
U_F7613: entity F port map(lamdaA => P(7)(613),lamdaB => P(7)(621),lamdaOut => P(6)(613));
U_F7614: entity F port map(lamdaA => P(7)(614),lamdaB => P(7)(622),lamdaOut => P(6)(614));
U_F7615: entity F port map(lamdaA => P(7)(615),lamdaB => P(7)(623),lamdaOut => P(6)(615));
U_G7616: entity G port map(lamdaA => P(7)(608),lamdaB => P(7)(616),s => s(7)(304),lamdaOut => P(6)(616));
U_G7617: entity G port map(lamdaA => P(7)(609),lamdaB => P(7)(617),s => s(7)(305),lamdaOut => P(6)(617));
U_G7618: entity G port map(lamdaA => P(7)(610),lamdaB => P(7)(618),s => s(7)(306),lamdaOut => P(6)(618));
U_G7619: entity G port map(lamdaA => P(7)(611),lamdaB => P(7)(619),s => s(7)(307),lamdaOut => P(6)(619));
U_G7620: entity G port map(lamdaA => P(7)(612),lamdaB => P(7)(620),s => s(7)(308),lamdaOut => P(6)(620));
U_G7621: entity G port map(lamdaA => P(7)(613),lamdaB => P(7)(621),s => s(7)(309),lamdaOut => P(6)(621));
U_G7622: entity G port map(lamdaA => P(7)(614),lamdaB => P(7)(622),s => s(7)(310),lamdaOut => P(6)(622));
U_G7623: entity G port map(lamdaA => P(7)(615),lamdaB => P(7)(623),s => s(7)(311),lamdaOut => P(6)(623));
U_F7624: entity F port map(lamdaA => P(7)(624),lamdaB => P(7)(632),lamdaOut => P(6)(624));
U_F7625: entity F port map(lamdaA => P(7)(625),lamdaB => P(7)(633),lamdaOut => P(6)(625));
U_F7626: entity F port map(lamdaA => P(7)(626),lamdaB => P(7)(634),lamdaOut => P(6)(626));
U_F7627: entity F port map(lamdaA => P(7)(627),lamdaB => P(7)(635),lamdaOut => P(6)(627));
U_F7628: entity F port map(lamdaA => P(7)(628),lamdaB => P(7)(636),lamdaOut => P(6)(628));
U_F7629: entity F port map(lamdaA => P(7)(629),lamdaB => P(7)(637),lamdaOut => P(6)(629));
U_F7630: entity F port map(lamdaA => P(7)(630),lamdaB => P(7)(638),lamdaOut => P(6)(630));
U_F7631: entity F port map(lamdaA => P(7)(631),lamdaB => P(7)(639),lamdaOut => P(6)(631));
U_G7632: entity G port map(lamdaA => P(7)(624),lamdaB => P(7)(632),s => s(7)(312),lamdaOut => P(6)(632));
U_G7633: entity G port map(lamdaA => P(7)(625),lamdaB => P(7)(633),s => s(7)(313),lamdaOut => P(6)(633));
U_G7634: entity G port map(lamdaA => P(7)(626),lamdaB => P(7)(634),s => s(7)(314),lamdaOut => P(6)(634));
U_G7635: entity G port map(lamdaA => P(7)(627),lamdaB => P(7)(635),s => s(7)(315),lamdaOut => P(6)(635));
U_G7636: entity G port map(lamdaA => P(7)(628),lamdaB => P(7)(636),s => s(7)(316),lamdaOut => P(6)(636));
U_G7637: entity G port map(lamdaA => P(7)(629),lamdaB => P(7)(637),s => s(7)(317),lamdaOut => P(6)(637));
U_G7638: entity G port map(lamdaA => P(7)(630),lamdaB => P(7)(638),s => s(7)(318),lamdaOut => P(6)(638));
U_G7639: entity G port map(lamdaA => P(7)(631),lamdaB => P(7)(639),s => s(7)(319),lamdaOut => P(6)(639));
U_F7640: entity F port map(lamdaA => P(7)(640),lamdaB => P(7)(648),lamdaOut => P(6)(640));
U_F7641: entity F port map(lamdaA => P(7)(641),lamdaB => P(7)(649),lamdaOut => P(6)(641));
U_F7642: entity F port map(lamdaA => P(7)(642),lamdaB => P(7)(650),lamdaOut => P(6)(642));
U_F7643: entity F port map(lamdaA => P(7)(643),lamdaB => P(7)(651),lamdaOut => P(6)(643));
U_F7644: entity F port map(lamdaA => P(7)(644),lamdaB => P(7)(652),lamdaOut => P(6)(644));
U_F7645: entity F port map(lamdaA => P(7)(645),lamdaB => P(7)(653),lamdaOut => P(6)(645));
U_F7646: entity F port map(lamdaA => P(7)(646),lamdaB => P(7)(654),lamdaOut => P(6)(646));
U_F7647: entity F port map(lamdaA => P(7)(647),lamdaB => P(7)(655),lamdaOut => P(6)(647));
U_G7648: entity G port map(lamdaA => P(7)(640),lamdaB => P(7)(648),s => s(7)(320),lamdaOut => P(6)(648));
U_G7649: entity G port map(lamdaA => P(7)(641),lamdaB => P(7)(649),s => s(7)(321),lamdaOut => P(6)(649));
U_G7650: entity G port map(lamdaA => P(7)(642),lamdaB => P(7)(650),s => s(7)(322),lamdaOut => P(6)(650));
U_G7651: entity G port map(lamdaA => P(7)(643),lamdaB => P(7)(651),s => s(7)(323),lamdaOut => P(6)(651));
U_G7652: entity G port map(lamdaA => P(7)(644),lamdaB => P(7)(652),s => s(7)(324),lamdaOut => P(6)(652));
U_G7653: entity G port map(lamdaA => P(7)(645),lamdaB => P(7)(653),s => s(7)(325),lamdaOut => P(6)(653));
U_G7654: entity G port map(lamdaA => P(7)(646),lamdaB => P(7)(654),s => s(7)(326),lamdaOut => P(6)(654));
U_G7655: entity G port map(lamdaA => P(7)(647),lamdaB => P(7)(655),s => s(7)(327),lamdaOut => P(6)(655));
U_F7656: entity F port map(lamdaA => P(7)(656),lamdaB => P(7)(664),lamdaOut => P(6)(656));
U_F7657: entity F port map(lamdaA => P(7)(657),lamdaB => P(7)(665),lamdaOut => P(6)(657));
U_F7658: entity F port map(lamdaA => P(7)(658),lamdaB => P(7)(666),lamdaOut => P(6)(658));
U_F7659: entity F port map(lamdaA => P(7)(659),lamdaB => P(7)(667),lamdaOut => P(6)(659));
U_F7660: entity F port map(lamdaA => P(7)(660),lamdaB => P(7)(668),lamdaOut => P(6)(660));
U_F7661: entity F port map(lamdaA => P(7)(661),lamdaB => P(7)(669),lamdaOut => P(6)(661));
U_F7662: entity F port map(lamdaA => P(7)(662),lamdaB => P(7)(670),lamdaOut => P(6)(662));
U_F7663: entity F port map(lamdaA => P(7)(663),lamdaB => P(7)(671),lamdaOut => P(6)(663));
U_G7664: entity G port map(lamdaA => P(7)(656),lamdaB => P(7)(664),s => s(7)(328),lamdaOut => P(6)(664));
U_G7665: entity G port map(lamdaA => P(7)(657),lamdaB => P(7)(665),s => s(7)(329),lamdaOut => P(6)(665));
U_G7666: entity G port map(lamdaA => P(7)(658),lamdaB => P(7)(666),s => s(7)(330),lamdaOut => P(6)(666));
U_G7667: entity G port map(lamdaA => P(7)(659),lamdaB => P(7)(667),s => s(7)(331),lamdaOut => P(6)(667));
U_G7668: entity G port map(lamdaA => P(7)(660),lamdaB => P(7)(668),s => s(7)(332),lamdaOut => P(6)(668));
U_G7669: entity G port map(lamdaA => P(7)(661),lamdaB => P(7)(669),s => s(7)(333),lamdaOut => P(6)(669));
U_G7670: entity G port map(lamdaA => P(7)(662),lamdaB => P(7)(670),s => s(7)(334),lamdaOut => P(6)(670));
U_G7671: entity G port map(lamdaA => P(7)(663),lamdaB => P(7)(671),s => s(7)(335),lamdaOut => P(6)(671));
U_F7672: entity F port map(lamdaA => P(7)(672),lamdaB => P(7)(680),lamdaOut => P(6)(672));
U_F7673: entity F port map(lamdaA => P(7)(673),lamdaB => P(7)(681),lamdaOut => P(6)(673));
U_F7674: entity F port map(lamdaA => P(7)(674),lamdaB => P(7)(682),lamdaOut => P(6)(674));
U_F7675: entity F port map(lamdaA => P(7)(675),lamdaB => P(7)(683),lamdaOut => P(6)(675));
U_F7676: entity F port map(lamdaA => P(7)(676),lamdaB => P(7)(684),lamdaOut => P(6)(676));
U_F7677: entity F port map(lamdaA => P(7)(677),lamdaB => P(7)(685),lamdaOut => P(6)(677));
U_F7678: entity F port map(lamdaA => P(7)(678),lamdaB => P(7)(686),lamdaOut => P(6)(678));
U_F7679: entity F port map(lamdaA => P(7)(679),lamdaB => P(7)(687),lamdaOut => P(6)(679));
U_G7680: entity G port map(lamdaA => P(7)(672),lamdaB => P(7)(680),s => s(7)(336),lamdaOut => P(6)(680));
U_G7681: entity G port map(lamdaA => P(7)(673),lamdaB => P(7)(681),s => s(7)(337),lamdaOut => P(6)(681));
U_G7682: entity G port map(lamdaA => P(7)(674),lamdaB => P(7)(682),s => s(7)(338),lamdaOut => P(6)(682));
U_G7683: entity G port map(lamdaA => P(7)(675),lamdaB => P(7)(683),s => s(7)(339),lamdaOut => P(6)(683));
U_G7684: entity G port map(lamdaA => P(7)(676),lamdaB => P(7)(684),s => s(7)(340),lamdaOut => P(6)(684));
U_G7685: entity G port map(lamdaA => P(7)(677),lamdaB => P(7)(685),s => s(7)(341),lamdaOut => P(6)(685));
U_G7686: entity G port map(lamdaA => P(7)(678),lamdaB => P(7)(686),s => s(7)(342),lamdaOut => P(6)(686));
U_G7687: entity G port map(lamdaA => P(7)(679),lamdaB => P(7)(687),s => s(7)(343),lamdaOut => P(6)(687));
U_F7688: entity F port map(lamdaA => P(7)(688),lamdaB => P(7)(696),lamdaOut => P(6)(688));
U_F7689: entity F port map(lamdaA => P(7)(689),lamdaB => P(7)(697),lamdaOut => P(6)(689));
U_F7690: entity F port map(lamdaA => P(7)(690),lamdaB => P(7)(698),lamdaOut => P(6)(690));
U_F7691: entity F port map(lamdaA => P(7)(691),lamdaB => P(7)(699),lamdaOut => P(6)(691));
U_F7692: entity F port map(lamdaA => P(7)(692),lamdaB => P(7)(700),lamdaOut => P(6)(692));
U_F7693: entity F port map(lamdaA => P(7)(693),lamdaB => P(7)(701),lamdaOut => P(6)(693));
U_F7694: entity F port map(lamdaA => P(7)(694),lamdaB => P(7)(702),lamdaOut => P(6)(694));
U_F7695: entity F port map(lamdaA => P(7)(695),lamdaB => P(7)(703),lamdaOut => P(6)(695));
U_G7696: entity G port map(lamdaA => P(7)(688),lamdaB => P(7)(696),s => s(7)(344),lamdaOut => P(6)(696));
U_G7697: entity G port map(lamdaA => P(7)(689),lamdaB => P(7)(697),s => s(7)(345),lamdaOut => P(6)(697));
U_G7698: entity G port map(lamdaA => P(7)(690),lamdaB => P(7)(698),s => s(7)(346),lamdaOut => P(6)(698));
U_G7699: entity G port map(lamdaA => P(7)(691),lamdaB => P(7)(699),s => s(7)(347),lamdaOut => P(6)(699));
U_G7700: entity G port map(lamdaA => P(7)(692),lamdaB => P(7)(700),s => s(7)(348),lamdaOut => P(6)(700));
U_G7701: entity G port map(lamdaA => P(7)(693),lamdaB => P(7)(701),s => s(7)(349),lamdaOut => P(6)(701));
U_G7702: entity G port map(lamdaA => P(7)(694),lamdaB => P(7)(702),s => s(7)(350),lamdaOut => P(6)(702));
U_G7703: entity G port map(lamdaA => P(7)(695),lamdaB => P(7)(703),s => s(7)(351),lamdaOut => P(6)(703));
U_F7704: entity F port map(lamdaA => P(7)(704),lamdaB => P(7)(712),lamdaOut => P(6)(704));
U_F7705: entity F port map(lamdaA => P(7)(705),lamdaB => P(7)(713),lamdaOut => P(6)(705));
U_F7706: entity F port map(lamdaA => P(7)(706),lamdaB => P(7)(714),lamdaOut => P(6)(706));
U_F7707: entity F port map(lamdaA => P(7)(707),lamdaB => P(7)(715),lamdaOut => P(6)(707));
U_F7708: entity F port map(lamdaA => P(7)(708),lamdaB => P(7)(716),lamdaOut => P(6)(708));
U_F7709: entity F port map(lamdaA => P(7)(709),lamdaB => P(7)(717),lamdaOut => P(6)(709));
U_F7710: entity F port map(lamdaA => P(7)(710),lamdaB => P(7)(718),lamdaOut => P(6)(710));
U_F7711: entity F port map(lamdaA => P(7)(711),lamdaB => P(7)(719),lamdaOut => P(6)(711));
U_G7712: entity G port map(lamdaA => P(7)(704),lamdaB => P(7)(712),s => s(7)(352),lamdaOut => P(6)(712));
U_G7713: entity G port map(lamdaA => P(7)(705),lamdaB => P(7)(713),s => s(7)(353),lamdaOut => P(6)(713));
U_G7714: entity G port map(lamdaA => P(7)(706),lamdaB => P(7)(714),s => s(7)(354),lamdaOut => P(6)(714));
U_G7715: entity G port map(lamdaA => P(7)(707),lamdaB => P(7)(715),s => s(7)(355),lamdaOut => P(6)(715));
U_G7716: entity G port map(lamdaA => P(7)(708),lamdaB => P(7)(716),s => s(7)(356),lamdaOut => P(6)(716));
U_G7717: entity G port map(lamdaA => P(7)(709),lamdaB => P(7)(717),s => s(7)(357),lamdaOut => P(6)(717));
U_G7718: entity G port map(lamdaA => P(7)(710),lamdaB => P(7)(718),s => s(7)(358),lamdaOut => P(6)(718));
U_G7719: entity G port map(lamdaA => P(7)(711),lamdaB => P(7)(719),s => s(7)(359),lamdaOut => P(6)(719));
U_F7720: entity F port map(lamdaA => P(7)(720),lamdaB => P(7)(728),lamdaOut => P(6)(720));
U_F7721: entity F port map(lamdaA => P(7)(721),lamdaB => P(7)(729),lamdaOut => P(6)(721));
U_F7722: entity F port map(lamdaA => P(7)(722),lamdaB => P(7)(730),lamdaOut => P(6)(722));
U_F7723: entity F port map(lamdaA => P(7)(723),lamdaB => P(7)(731),lamdaOut => P(6)(723));
U_F7724: entity F port map(lamdaA => P(7)(724),lamdaB => P(7)(732),lamdaOut => P(6)(724));
U_F7725: entity F port map(lamdaA => P(7)(725),lamdaB => P(7)(733),lamdaOut => P(6)(725));
U_F7726: entity F port map(lamdaA => P(7)(726),lamdaB => P(7)(734),lamdaOut => P(6)(726));
U_F7727: entity F port map(lamdaA => P(7)(727),lamdaB => P(7)(735),lamdaOut => P(6)(727));
U_G7728: entity G port map(lamdaA => P(7)(720),lamdaB => P(7)(728),s => s(7)(360),lamdaOut => P(6)(728));
U_G7729: entity G port map(lamdaA => P(7)(721),lamdaB => P(7)(729),s => s(7)(361),lamdaOut => P(6)(729));
U_G7730: entity G port map(lamdaA => P(7)(722),lamdaB => P(7)(730),s => s(7)(362),lamdaOut => P(6)(730));
U_G7731: entity G port map(lamdaA => P(7)(723),lamdaB => P(7)(731),s => s(7)(363),lamdaOut => P(6)(731));
U_G7732: entity G port map(lamdaA => P(7)(724),lamdaB => P(7)(732),s => s(7)(364),lamdaOut => P(6)(732));
U_G7733: entity G port map(lamdaA => P(7)(725),lamdaB => P(7)(733),s => s(7)(365),lamdaOut => P(6)(733));
U_G7734: entity G port map(lamdaA => P(7)(726),lamdaB => P(7)(734),s => s(7)(366),lamdaOut => P(6)(734));
U_G7735: entity G port map(lamdaA => P(7)(727),lamdaB => P(7)(735),s => s(7)(367),lamdaOut => P(6)(735));
U_F7736: entity F port map(lamdaA => P(7)(736),lamdaB => P(7)(744),lamdaOut => P(6)(736));
U_F7737: entity F port map(lamdaA => P(7)(737),lamdaB => P(7)(745),lamdaOut => P(6)(737));
U_F7738: entity F port map(lamdaA => P(7)(738),lamdaB => P(7)(746),lamdaOut => P(6)(738));
U_F7739: entity F port map(lamdaA => P(7)(739),lamdaB => P(7)(747),lamdaOut => P(6)(739));
U_F7740: entity F port map(lamdaA => P(7)(740),lamdaB => P(7)(748),lamdaOut => P(6)(740));
U_F7741: entity F port map(lamdaA => P(7)(741),lamdaB => P(7)(749),lamdaOut => P(6)(741));
U_F7742: entity F port map(lamdaA => P(7)(742),lamdaB => P(7)(750),lamdaOut => P(6)(742));
U_F7743: entity F port map(lamdaA => P(7)(743),lamdaB => P(7)(751),lamdaOut => P(6)(743));
U_G7744: entity G port map(lamdaA => P(7)(736),lamdaB => P(7)(744),s => s(7)(368),lamdaOut => P(6)(744));
U_G7745: entity G port map(lamdaA => P(7)(737),lamdaB => P(7)(745),s => s(7)(369),lamdaOut => P(6)(745));
U_G7746: entity G port map(lamdaA => P(7)(738),lamdaB => P(7)(746),s => s(7)(370),lamdaOut => P(6)(746));
U_G7747: entity G port map(lamdaA => P(7)(739),lamdaB => P(7)(747),s => s(7)(371),lamdaOut => P(6)(747));
U_G7748: entity G port map(lamdaA => P(7)(740),lamdaB => P(7)(748),s => s(7)(372),lamdaOut => P(6)(748));
U_G7749: entity G port map(lamdaA => P(7)(741),lamdaB => P(7)(749),s => s(7)(373),lamdaOut => P(6)(749));
U_G7750: entity G port map(lamdaA => P(7)(742),lamdaB => P(7)(750),s => s(7)(374),lamdaOut => P(6)(750));
U_G7751: entity G port map(lamdaA => P(7)(743),lamdaB => P(7)(751),s => s(7)(375),lamdaOut => P(6)(751));
U_F7752: entity F port map(lamdaA => P(7)(752),lamdaB => P(7)(760),lamdaOut => P(6)(752));
U_F7753: entity F port map(lamdaA => P(7)(753),lamdaB => P(7)(761),lamdaOut => P(6)(753));
U_F7754: entity F port map(lamdaA => P(7)(754),lamdaB => P(7)(762),lamdaOut => P(6)(754));
U_F7755: entity F port map(lamdaA => P(7)(755),lamdaB => P(7)(763),lamdaOut => P(6)(755));
U_F7756: entity F port map(lamdaA => P(7)(756),lamdaB => P(7)(764),lamdaOut => P(6)(756));
U_F7757: entity F port map(lamdaA => P(7)(757),lamdaB => P(7)(765),lamdaOut => P(6)(757));
U_F7758: entity F port map(lamdaA => P(7)(758),lamdaB => P(7)(766),lamdaOut => P(6)(758));
U_F7759: entity F port map(lamdaA => P(7)(759),lamdaB => P(7)(767),lamdaOut => P(6)(759));
U_G7760: entity G port map(lamdaA => P(7)(752),lamdaB => P(7)(760),s => s(7)(376),lamdaOut => P(6)(760));
U_G7761: entity G port map(lamdaA => P(7)(753),lamdaB => P(7)(761),s => s(7)(377),lamdaOut => P(6)(761));
U_G7762: entity G port map(lamdaA => P(7)(754),lamdaB => P(7)(762),s => s(7)(378),lamdaOut => P(6)(762));
U_G7763: entity G port map(lamdaA => P(7)(755),lamdaB => P(7)(763),s => s(7)(379),lamdaOut => P(6)(763));
U_G7764: entity G port map(lamdaA => P(7)(756),lamdaB => P(7)(764),s => s(7)(380),lamdaOut => P(6)(764));
U_G7765: entity G port map(lamdaA => P(7)(757),lamdaB => P(7)(765),s => s(7)(381),lamdaOut => P(6)(765));
U_G7766: entity G port map(lamdaA => P(7)(758),lamdaB => P(7)(766),s => s(7)(382),lamdaOut => P(6)(766));
U_G7767: entity G port map(lamdaA => P(7)(759),lamdaB => P(7)(767),s => s(7)(383),lamdaOut => P(6)(767));
U_F7768: entity F port map(lamdaA => P(7)(768),lamdaB => P(7)(776),lamdaOut => P(6)(768));
U_F7769: entity F port map(lamdaA => P(7)(769),lamdaB => P(7)(777),lamdaOut => P(6)(769));
U_F7770: entity F port map(lamdaA => P(7)(770),lamdaB => P(7)(778),lamdaOut => P(6)(770));
U_F7771: entity F port map(lamdaA => P(7)(771),lamdaB => P(7)(779),lamdaOut => P(6)(771));
U_F7772: entity F port map(lamdaA => P(7)(772),lamdaB => P(7)(780),lamdaOut => P(6)(772));
U_F7773: entity F port map(lamdaA => P(7)(773),lamdaB => P(7)(781),lamdaOut => P(6)(773));
U_F7774: entity F port map(lamdaA => P(7)(774),lamdaB => P(7)(782),lamdaOut => P(6)(774));
U_F7775: entity F port map(lamdaA => P(7)(775),lamdaB => P(7)(783),lamdaOut => P(6)(775));
U_G7776: entity G port map(lamdaA => P(7)(768),lamdaB => P(7)(776),s => s(7)(384),lamdaOut => P(6)(776));
U_G7777: entity G port map(lamdaA => P(7)(769),lamdaB => P(7)(777),s => s(7)(385),lamdaOut => P(6)(777));
U_G7778: entity G port map(lamdaA => P(7)(770),lamdaB => P(7)(778),s => s(7)(386),lamdaOut => P(6)(778));
U_G7779: entity G port map(lamdaA => P(7)(771),lamdaB => P(7)(779),s => s(7)(387),lamdaOut => P(6)(779));
U_G7780: entity G port map(lamdaA => P(7)(772),lamdaB => P(7)(780),s => s(7)(388),lamdaOut => P(6)(780));
U_G7781: entity G port map(lamdaA => P(7)(773),lamdaB => P(7)(781),s => s(7)(389),lamdaOut => P(6)(781));
U_G7782: entity G port map(lamdaA => P(7)(774),lamdaB => P(7)(782),s => s(7)(390),lamdaOut => P(6)(782));
U_G7783: entity G port map(lamdaA => P(7)(775),lamdaB => P(7)(783),s => s(7)(391),lamdaOut => P(6)(783));
U_F7784: entity F port map(lamdaA => P(7)(784),lamdaB => P(7)(792),lamdaOut => P(6)(784));
U_F7785: entity F port map(lamdaA => P(7)(785),lamdaB => P(7)(793),lamdaOut => P(6)(785));
U_F7786: entity F port map(lamdaA => P(7)(786),lamdaB => P(7)(794),lamdaOut => P(6)(786));
U_F7787: entity F port map(lamdaA => P(7)(787),lamdaB => P(7)(795),lamdaOut => P(6)(787));
U_F7788: entity F port map(lamdaA => P(7)(788),lamdaB => P(7)(796),lamdaOut => P(6)(788));
U_F7789: entity F port map(lamdaA => P(7)(789),lamdaB => P(7)(797),lamdaOut => P(6)(789));
U_F7790: entity F port map(lamdaA => P(7)(790),lamdaB => P(7)(798),lamdaOut => P(6)(790));
U_F7791: entity F port map(lamdaA => P(7)(791),lamdaB => P(7)(799),lamdaOut => P(6)(791));
U_G7792: entity G port map(lamdaA => P(7)(784),lamdaB => P(7)(792),s => s(7)(392),lamdaOut => P(6)(792));
U_G7793: entity G port map(lamdaA => P(7)(785),lamdaB => P(7)(793),s => s(7)(393),lamdaOut => P(6)(793));
U_G7794: entity G port map(lamdaA => P(7)(786),lamdaB => P(7)(794),s => s(7)(394),lamdaOut => P(6)(794));
U_G7795: entity G port map(lamdaA => P(7)(787),lamdaB => P(7)(795),s => s(7)(395),lamdaOut => P(6)(795));
U_G7796: entity G port map(lamdaA => P(7)(788),lamdaB => P(7)(796),s => s(7)(396),lamdaOut => P(6)(796));
U_G7797: entity G port map(lamdaA => P(7)(789),lamdaB => P(7)(797),s => s(7)(397),lamdaOut => P(6)(797));
U_G7798: entity G port map(lamdaA => P(7)(790),lamdaB => P(7)(798),s => s(7)(398),lamdaOut => P(6)(798));
U_G7799: entity G port map(lamdaA => P(7)(791),lamdaB => P(7)(799),s => s(7)(399),lamdaOut => P(6)(799));
U_F7800: entity F port map(lamdaA => P(7)(800),lamdaB => P(7)(808),lamdaOut => P(6)(800));
U_F7801: entity F port map(lamdaA => P(7)(801),lamdaB => P(7)(809),lamdaOut => P(6)(801));
U_F7802: entity F port map(lamdaA => P(7)(802),lamdaB => P(7)(810),lamdaOut => P(6)(802));
U_F7803: entity F port map(lamdaA => P(7)(803),lamdaB => P(7)(811),lamdaOut => P(6)(803));
U_F7804: entity F port map(lamdaA => P(7)(804),lamdaB => P(7)(812),lamdaOut => P(6)(804));
U_F7805: entity F port map(lamdaA => P(7)(805),lamdaB => P(7)(813),lamdaOut => P(6)(805));
U_F7806: entity F port map(lamdaA => P(7)(806),lamdaB => P(7)(814),lamdaOut => P(6)(806));
U_F7807: entity F port map(lamdaA => P(7)(807),lamdaB => P(7)(815),lamdaOut => P(6)(807));
U_G7808: entity G port map(lamdaA => P(7)(800),lamdaB => P(7)(808),s => s(7)(400),lamdaOut => P(6)(808));
U_G7809: entity G port map(lamdaA => P(7)(801),lamdaB => P(7)(809),s => s(7)(401),lamdaOut => P(6)(809));
U_G7810: entity G port map(lamdaA => P(7)(802),lamdaB => P(7)(810),s => s(7)(402),lamdaOut => P(6)(810));
U_G7811: entity G port map(lamdaA => P(7)(803),lamdaB => P(7)(811),s => s(7)(403),lamdaOut => P(6)(811));
U_G7812: entity G port map(lamdaA => P(7)(804),lamdaB => P(7)(812),s => s(7)(404),lamdaOut => P(6)(812));
U_G7813: entity G port map(lamdaA => P(7)(805),lamdaB => P(7)(813),s => s(7)(405),lamdaOut => P(6)(813));
U_G7814: entity G port map(lamdaA => P(7)(806),lamdaB => P(7)(814),s => s(7)(406),lamdaOut => P(6)(814));
U_G7815: entity G port map(lamdaA => P(7)(807),lamdaB => P(7)(815),s => s(7)(407),lamdaOut => P(6)(815));
U_F7816: entity F port map(lamdaA => P(7)(816),lamdaB => P(7)(824),lamdaOut => P(6)(816));
U_F7817: entity F port map(lamdaA => P(7)(817),lamdaB => P(7)(825),lamdaOut => P(6)(817));
U_F7818: entity F port map(lamdaA => P(7)(818),lamdaB => P(7)(826),lamdaOut => P(6)(818));
U_F7819: entity F port map(lamdaA => P(7)(819),lamdaB => P(7)(827),lamdaOut => P(6)(819));
U_F7820: entity F port map(lamdaA => P(7)(820),lamdaB => P(7)(828),lamdaOut => P(6)(820));
U_F7821: entity F port map(lamdaA => P(7)(821),lamdaB => P(7)(829),lamdaOut => P(6)(821));
U_F7822: entity F port map(lamdaA => P(7)(822),lamdaB => P(7)(830),lamdaOut => P(6)(822));
U_F7823: entity F port map(lamdaA => P(7)(823),lamdaB => P(7)(831),lamdaOut => P(6)(823));
U_G7824: entity G port map(lamdaA => P(7)(816),lamdaB => P(7)(824),s => s(7)(408),lamdaOut => P(6)(824));
U_G7825: entity G port map(lamdaA => P(7)(817),lamdaB => P(7)(825),s => s(7)(409),lamdaOut => P(6)(825));
U_G7826: entity G port map(lamdaA => P(7)(818),lamdaB => P(7)(826),s => s(7)(410),lamdaOut => P(6)(826));
U_G7827: entity G port map(lamdaA => P(7)(819),lamdaB => P(7)(827),s => s(7)(411),lamdaOut => P(6)(827));
U_G7828: entity G port map(lamdaA => P(7)(820),lamdaB => P(7)(828),s => s(7)(412),lamdaOut => P(6)(828));
U_G7829: entity G port map(lamdaA => P(7)(821),lamdaB => P(7)(829),s => s(7)(413),lamdaOut => P(6)(829));
U_G7830: entity G port map(lamdaA => P(7)(822),lamdaB => P(7)(830),s => s(7)(414),lamdaOut => P(6)(830));
U_G7831: entity G port map(lamdaA => P(7)(823),lamdaB => P(7)(831),s => s(7)(415),lamdaOut => P(6)(831));
U_F7832: entity F port map(lamdaA => P(7)(832),lamdaB => P(7)(840),lamdaOut => P(6)(832));
U_F7833: entity F port map(lamdaA => P(7)(833),lamdaB => P(7)(841),lamdaOut => P(6)(833));
U_F7834: entity F port map(lamdaA => P(7)(834),lamdaB => P(7)(842),lamdaOut => P(6)(834));
U_F7835: entity F port map(lamdaA => P(7)(835),lamdaB => P(7)(843),lamdaOut => P(6)(835));
U_F7836: entity F port map(lamdaA => P(7)(836),lamdaB => P(7)(844),lamdaOut => P(6)(836));
U_F7837: entity F port map(lamdaA => P(7)(837),lamdaB => P(7)(845),lamdaOut => P(6)(837));
U_F7838: entity F port map(lamdaA => P(7)(838),lamdaB => P(7)(846),lamdaOut => P(6)(838));
U_F7839: entity F port map(lamdaA => P(7)(839),lamdaB => P(7)(847),lamdaOut => P(6)(839));
U_G7840: entity G port map(lamdaA => P(7)(832),lamdaB => P(7)(840),s => s(7)(416),lamdaOut => P(6)(840));
U_G7841: entity G port map(lamdaA => P(7)(833),lamdaB => P(7)(841),s => s(7)(417),lamdaOut => P(6)(841));
U_G7842: entity G port map(lamdaA => P(7)(834),lamdaB => P(7)(842),s => s(7)(418),lamdaOut => P(6)(842));
U_G7843: entity G port map(lamdaA => P(7)(835),lamdaB => P(7)(843),s => s(7)(419),lamdaOut => P(6)(843));
U_G7844: entity G port map(lamdaA => P(7)(836),lamdaB => P(7)(844),s => s(7)(420),lamdaOut => P(6)(844));
U_G7845: entity G port map(lamdaA => P(7)(837),lamdaB => P(7)(845),s => s(7)(421),lamdaOut => P(6)(845));
U_G7846: entity G port map(lamdaA => P(7)(838),lamdaB => P(7)(846),s => s(7)(422),lamdaOut => P(6)(846));
U_G7847: entity G port map(lamdaA => P(7)(839),lamdaB => P(7)(847),s => s(7)(423),lamdaOut => P(6)(847));
U_F7848: entity F port map(lamdaA => P(7)(848),lamdaB => P(7)(856),lamdaOut => P(6)(848));
U_F7849: entity F port map(lamdaA => P(7)(849),lamdaB => P(7)(857),lamdaOut => P(6)(849));
U_F7850: entity F port map(lamdaA => P(7)(850),lamdaB => P(7)(858),lamdaOut => P(6)(850));
U_F7851: entity F port map(lamdaA => P(7)(851),lamdaB => P(7)(859),lamdaOut => P(6)(851));
U_F7852: entity F port map(lamdaA => P(7)(852),lamdaB => P(7)(860),lamdaOut => P(6)(852));
U_F7853: entity F port map(lamdaA => P(7)(853),lamdaB => P(7)(861),lamdaOut => P(6)(853));
U_F7854: entity F port map(lamdaA => P(7)(854),lamdaB => P(7)(862),lamdaOut => P(6)(854));
U_F7855: entity F port map(lamdaA => P(7)(855),lamdaB => P(7)(863),lamdaOut => P(6)(855));
U_G7856: entity G port map(lamdaA => P(7)(848),lamdaB => P(7)(856),s => s(7)(424),lamdaOut => P(6)(856));
U_G7857: entity G port map(lamdaA => P(7)(849),lamdaB => P(7)(857),s => s(7)(425),lamdaOut => P(6)(857));
U_G7858: entity G port map(lamdaA => P(7)(850),lamdaB => P(7)(858),s => s(7)(426),lamdaOut => P(6)(858));
U_G7859: entity G port map(lamdaA => P(7)(851),lamdaB => P(7)(859),s => s(7)(427),lamdaOut => P(6)(859));
U_G7860: entity G port map(lamdaA => P(7)(852),lamdaB => P(7)(860),s => s(7)(428),lamdaOut => P(6)(860));
U_G7861: entity G port map(lamdaA => P(7)(853),lamdaB => P(7)(861),s => s(7)(429),lamdaOut => P(6)(861));
U_G7862: entity G port map(lamdaA => P(7)(854),lamdaB => P(7)(862),s => s(7)(430),lamdaOut => P(6)(862));
U_G7863: entity G port map(lamdaA => P(7)(855),lamdaB => P(7)(863),s => s(7)(431),lamdaOut => P(6)(863));
U_F7864: entity F port map(lamdaA => P(7)(864),lamdaB => P(7)(872),lamdaOut => P(6)(864));
U_F7865: entity F port map(lamdaA => P(7)(865),lamdaB => P(7)(873),lamdaOut => P(6)(865));
U_F7866: entity F port map(lamdaA => P(7)(866),lamdaB => P(7)(874),lamdaOut => P(6)(866));
U_F7867: entity F port map(lamdaA => P(7)(867),lamdaB => P(7)(875),lamdaOut => P(6)(867));
U_F7868: entity F port map(lamdaA => P(7)(868),lamdaB => P(7)(876),lamdaOut => P(6)(868));
U_F7869: entity F port map(lamdaA => P(7)(869),lamdaB => P(7)(877),lamdaOut => P(6)(869));
U_F7870: entity F port map(lamdaA => P(7)(870),lamdaB => P(7)(878),lamdaOut => P(6)(870));
U_F7871: entity F port map(lamdaA => P(7)(871),lamdaB => P(7)(879),lamdaOut => P(6)(871));
U_G7872: entity G port map(lamdaA => P(7)(864),lamdaB => P(7)(872),s => s(7)(432),lamdaOut => P(6)(872));
U_G7873: entity G port map(lamdaA => P(7)(865),lamdaB => P(7)(873),s => s(7)(433),lamdaOut => P(6)(873));
U_G7874: entity G port map(lamdaA => P(7)(866),lamdaB => P(7)(874),s => s(7)(434),lamdaOut => P(6)(874));
U_G7875: entity G port map(lamdaA => P(7)(867),lamdaB => P(7)(875),s => s(7)(435),lamdaOut => P(6)(875));
U_G7876: entity G port map(lamdaA => P(7)(868),lamdaB => P(7)(876),s => s(7)(436),lamdaOut => P(6)(876));
U_G7877: entity G port map(lamdaA => P(7)(869),lamdaB => P(7)(877),s => s(7)(437),lamdaOut => P(6)(877));
U_G7878: entity G port map(lamdaA => P(7)(870),lamdaB => P(7)(878),s => s(7)(438),lamdaOut => P(6)(878));
U_G7879: entity G port map(lamdaA => P(7)(871),lamdaB => P(7)(879),s => s(7)(439),lamdaOut => P(6)(879));
U_F7880: entity F port map(lamdaA => P(7)(880),lamdaB => P(7)(888),lamdaOut => P(6)(880));
U_F7881: entity F port map(lamdaA => P(7)(881),lamdaB => P(7)(889),lamdaOut => P(6)(881));
U_F7882: entity F port map(lamdaA => P(7)(882),lamdaB => P(7)(890),lamdaOut => P(6)(882));
U_F7883: entity F port map(lamdaA => P(7)(883),lamdaB => P(7)(891),lamdaOut => P(6)(883));
U_F7884: entity F port map(lamdaA => P(7)(884),lamdaB => P(7)(892),lamdaOut => P(6)(884));
U_F7885: entity F port map(lamdaA => P(7)(885),lamdaB => P(7)(893),lamdaOut => P(6)(885));
U_F7886: entity F port map(lamdaA => P(7)(886),lamdaB => P(7)(894),lamdaOut => P(6)(886));
U_F7887: entity F port map(lamdaA => P(7)(887),lamdaB => P(7)(895),lamdaOut => P(6)(887));
U_G7888: entity G port map(lamdaA => P(7)(880),lamdaB => P(7)(888),s => s(7)(440),lamdaOut => P(6)(888));
U_G7889: entity G port map(lamdaA => P(7)(881),lamdaB => P(7)(889),s => s(7)(441),lamdaOut => P(6)(889));
U_G7890: entity G port map(lamdaA => P(7)(882),lamdaB => P(7)(890),s => s(7)(442),lamdaOut => P(6)(890));
U_G7891: entity G port map(lamdaA => P(7)(883),lamdaB => P(7)(891),s => s(7)(443),lamdaOut => P(6)(891));
U_G7892: entity G port map(lamdaA => P(7)(884),lamdaB => P(7)(892),s => s(7)(444),lamdaOut => P(6)(892));
U_G7893: entity G port map(lamdaA => P(7)(885),lamdaB => P(7)(893),s => s(7)(445),lamdaOut => P(6)(893));
U_G7894: entity G port map(lamdaA => P(7)(886),lamdaB => P(7)(894),s => s(7)(446),lamdaOut => P(6)(894));
U_G7895: entity G port map(lamdaA => P(7)(887),lamdaB => P(7)(895),s => s(7)(447),lamdaOut => P(6)(895));
U_F7896: entity F port map(lamdaA => P(7)(896),lamdaB => P(7)(904),lamdaOut => P(6)(896));
U_F7897: entity F port map(lamdaA => P(7)(897),lamdaB => P(7)(905),lamdaOut => P(6)(897));
U_F7898: entity F port map(lamdaA => P(7)(898),lamdaB => P(7)(906),lamdaOut => P(6)(898));
U_F7899: entity F port map(lamdaA => P(7)(899),lamdaB => P(7)(907),lamdaOut => P(6)(899));
U_F7900: entity F port map(lamdaA => P(7)(900),lamdaB => P(7)(908),lamdaOut => P(6)(900));
U_F7901: entity F port map(lamdaA => P(7)(901),lamdaB => P(7)(909),lamdaOut => P(6)(901));
U_F7902: entity F port map(lamdaA => P(7)(902),lamdaB => P(7)(910),lamdaOut => P(6)(902));
U_F7903: entity F port map(lamdaA => P(7)(903),lamdaB => P(7)(911),lamdaOut => P(6)(903));
U_G7904: entity G port map(lamdaA => P(7)(896),lamdaB => P(7)(904),s => s(7)(448),lamdaOut => P(6)(904));
U_G7905: entity G port map(lamdaA => P(7)(897),lamdaB => P(7)(905),s => s(7)(449),lamdaOut => P(6)(905));
U_G7906: entity G port map(lamdaA => P(7)(898),lamdaB => P(7)(906),s => s(7)(450),lamdaOut => P(6)(906));
U_G7907: entity G port map(lamdaA => P(7)(899),lamdaB => P(7)(907),s => s(7)(451),lamdaOut => P(6)(907));
U_G7908: entity G port map(lamdaA => P(7)(900),lamdaB => P(7)(908),s => s(7)(452),lamdaOut => P(6)(908));
U_G7909: entity G port map(lamdaA => P(7)(901),lamdaB => P(7)(909),s => s(7)(453),lamdaOut => P(6)(909));
U_G7910: entity G port map(lamdaA => P(7)(902),lamdaB => P(7)(910),s => s(7)(454),lamdaOut => P(6)(910));
U_G7911: entity G port map(lamdaA => P(7)(903),lamdaB => P(7)(911),s => s(7)(455),lamdaOut => P(6)(911));
U_F7912: entity F port map(lamdaA => P(7)(912),lamdaB => P(7)(920),lamdaOut => P(6)(912));
U_F7913: entity F port map(lamdaA => P(7)(913),lamdaB => P(7)(921),lamdaOut => P(6)(913));
U_F7914: entity F port map(lamdaA => P(7)(914),lamdaB => P(7)(922),lamdaOut => P(6)(914));
U_F7915: entity F port map(lamdaA => P(7)(915),lamdaB => P(7)(923),lamdaOut => P(6)(915));
U_F7916: entity F port map(lamdaA => P(7)(916),lamdaB => P(7)(924),lamdaOut => P(6)(916));
U_F7917: entity F port map(lamdaA => P(7)(917),lamdaB => P(7)(925),lamdaOut => P(6)(917));
U_F7918: entity F port map(lamdaA => P(7)(918),lamdaB => P(7)(926),lamdaOut => P(6)(918));
U_F7919: entity F port map(lamdaA => P(7)(919),lamdaB => P(7)(927),lamdaOut => P(6)(919));
U_G7920: entity G port map(lamdaA => P(7)(912),lamdaB => P(7)(920),s => s(7)(456),lamdaOut => P(6)(920));
U_G7921: entity G port map(lamdaA => P(7)(913),lamdaB => P(7)(921),s => s(7)(457),lamdaOut => P(6)(921));
U_G7922: entity G port map(lamdaA => P(7)(914),lamdaB => P(7)(922),s => s(7)(458),lamdaOut => P(6)(922));
U_G7923: entity G port map(lamdaA => P(7)(915),lamdaB => P(7)(923),s => s(7)(459),lamdaOut => P(6)(923));
U_G7924: entity G port map(lamdaA => P(7)(916),lamdaB => P(7)(924),s => s(7)(460),lamdaOut => P(6)(924));
U_G7925: entity G port map(lamdaA => P(7)(917),lamdaB => P(7)(925),s => s(7)(461),lamdaOut => P(6)(925));
U_G7926: entity G port map(lamdaA => P(7)(918),lamdaB => P(7)(926),s => s(7)(462),lamdaOut => P(6)(926));
U_G7927: entity G port map(lamdaA => P(7)(919),lamdaB => P(7)(927),s => s(7)(463),lamdaOut => P(6)(927));
U_F7928: entity F port map(lamdaA => P(7)(928),lamdaB => P(7)(936),lamdaOut => P(6)(928));
U_F7929: entity F port map(lamdaA => P(7)(929),lamdaB => P(7)(937),lamdaOut => P(6)(929));
U_F7930: entity F port map(lamdaA => P(7)(930),lamdaB => P(7)(938),lamdaOut => P(6)(930));
U_F7931: entity F port map(lamdaA => P(7)(931),lamdaB => P(7)(939),lamdaOut => P(6)(931));
U_F7932: entity F port map(lamdaA => P(7)(932),lamdaB => P(7)(940),lamdaOut => P(6)(932));
U_F7933: entity F port map(lamdaA => P(7)(933),lamdaB => P(7)(941),lamdaOut => P(6)(933));
U_F7934: entity F port map(lamdaA => P(7)(934),lamdaB => P(7)(942),lamdaOut => P(6)(934));
U_F7935: entity F port map(lamdaA => P(7)(935),lamdaB => P(7)(943),lamdaOut => P(6)(935));
U_G7936: entity G port map(lamdaA => P(7)(928),lamdaB => P(7)(936),s => s(7)(464),lamdaOut => P(6)(936));
U_G7937: entity G port map(lamdaA => P(7)(929),lamdaB => P(7)(937),s => s(7)(465),lamdaOut => P(6)(937));
U_G7938: entity G port map(lamdaA => P(7)(930),lamdaB => P(7)(938),s => s(7)(466),lamdaOut => P(6)(938));
U_G7939: entity G port map(lamdaA => P(7)(931),lamdaB => P(7)(939),s => s(7)(467),lamdaOut => P(6)(939));
U_G7940: entity G port map(lamdaA => P(7)(932),lamdaB => P(7)(940),s => s(7)(468),lamdaOut => P(6)(940));
U_G7941: entity G port map(lamdaA => P(7)(933),lamdaB => P(7)(941),s => s(7)(469),lamdaOut => P(6)(941));
U_G7942: entity G port map(lamdaA => P(7)(934),lamdaB => P(7)(942),s => s(7)(470),lamdaOut => P(6)(942));
U_G7943: entity G port map(lamdaA => P(7)(935),lamdaB => P(7)(943),s => s(7)(471),lamdaOut => P(6)(943));
U_F7944: entity F port map(lamdaA => P(7)(944),lamdaB => P(7)(952),lamdaOut => P(6)(944));
U_F7945: entity F port map(lamdaA => P(7)(945),lamdaB => P(7)(953),lamdaOut => P(6)(945));
U_F7946: entity F port map(lamdaA => P(7)(946),lamdaB => P(7)(954),lamdaOut => P(6)(946));
U_F7947: entity F port map(lamdaA => P(7)(947),lamdaB => P(7)(955),lamdaOut => P(6)(947));
U_F7948: entity F port map(lamdaA => P(7)(948),lamdaB => P(7)(956),lamdaOut => P(6)(948));
U_F7949: entity F port map(lamdaA => P(7)(949),lamdaB => P(7)(957),lamdaOut => P(6)(949));
U_F7950: entity F port map(lamdaA => P(7)(950),lamdaB => P(7)(958),lamdaOut => P(6)(950));
U_F7951: entity F port map(lamdaA => P(7)(951),lamdaB => P(7)(959),lamdaOut => P(6)(951));
U_G7952: entity G port map(lamdaA => P(7)(944),lamdaB => P(7)(952),s => s(7)(472),lamdaOut => P(6)(952));
U_G7953: entity G port map(lamdaA => P(7)(945),lamdaB => P(7)(953),s => s(7)(473),lamdaOut => P(6)(953));
U_G7954: entity G port map(lamdaA => P(7)(946),lamdaB => P(7)(954),s => s(7)(474),lamdaOut => P(6)(954));
U_G7955: entity G port map(lamdaA => P(7)(947),lamdaB => P(7)(955),s => s(7)(475),lamdaOut => P(6)(955));
U_G7956: entity G port map(lamdaA => P(7)(948),lamdaB => P(7)(956),s => s(7)(476),lamdaOut => P(6)(956));
U_G7957: entity G port map(lamdaA => P(7)(949),lamdaB => P(7)(957),s => s(7)(477),lamdaOut => P(6)(957));
U_G7958: entity G port map(lamdaA => P(7)(950),lamdaB => P(7)(958),s => s(7)(478),lamdaOut => P(6)(958));
U_G7959: entity G port map(lamdaA => P(7)(951),lamdaB => P(7)(959),s => s(7)(479),lamdaOut => P(6)(959));
U_F7960: entity F port map(lamdaA => P(7)(960),lamdaB => P(7)(968),lamdaOut => P(6)(960));
U_F7961: entity F port map(lamdaA => P(7)(961),lamdaB => P(7)(969),lamdaOut => P(6)(961));
U_F7962: entity F port map(lamdaA => P(7)(962),lamdaB => P(7)(970),lamdaOut => P(6)(962));
U_F7963: entity F port map(lamdaA => P(7)(963),lamdaB => P(7)(971),lamdaOut => P(6)(963));
U_F7964: entity F port map(lamdaA => P(7)(964),lamdaB => P(7)(972),lamdaOut => P(6)(964));
U_F7965: entity F port map(lamdaA => P(7)(965),lamdaB => P(7)(973),lamdaOut => P(6)(965));
U_F7966: entity F port map(lamdaA => P(7)(966),lamdaB => P(7)(974),lamdaOut => P(6)(966));
U_F7967: entity F port map(lamdaA => P(7)(967),lamdaB => P(7)(975),lamdaOut => P(6)(967));
U_G7968: entity G port map(lamdaA => P(7)(960),lamdaB => P(7)(968),s => s(7)(480),lamdaOut => P(6)(968));
U_G7969: entity G port map(lamdaA => P(7)(961),lamdaB => P(7)(969),s => s(7)(481),lamdaOut => P(6)(969));
U_G7970: entity G port map(lamdaA => P(7)(962),lamdaB => P(7)(970),s => s(7)(482),lamdaOut => P(6)(970));
U_G7971: entity G port map(lamdaA => P(7)(963),lamdaB => P(7)(971),s => s(7)(483),lamdaOut => P(6)(971));
U_G7972: entity G port map(lamdaA => P(7)(964),lamdaB => P(7)(972),s => s(7)(484),lamdaOut => P(6)(972));
U_G7973: entity G port map(lamdaA => P(7)(965),lamdaB => P(7)(973),s => s(7)(485),lamdaOut => P(6)(973));
U_G7974: entity G port map(lamdaA => P(7)(966),lamdaB => P(7)(974),s => s(7)(486),lamdaOut => P(6)(974));
U_G7975: entity G port map(lamdaA => P(7)(967),lamdaB => P(7)(975),s => s(7)(487),lamdaOut => P(6)(975));
U_F7976: entity F port map(lamdaA => P(7)(976),lamdaB => P(7)(984),lamdaOut => P(6)(976));
U_F7977: entity F port map(lamdaA => P(7)(977),lamdaB => P(7)(985),lamdaOut => P(6)(977));
U_F7978: entity F port map(lamdaA => P(7)(978),lamdaB => P(7)(986),lamdaOut => P(6)(978));
U_F7979: entity F port map(lamdaA => P(7)(979),lamdaB => P(7)(987),lamdaOut => P(6)(979));
U_F7980: entity F port map(lamdaA => P(7)(980),lamdaB => P(7)(988),lamdaOut => P(6)(980));
U_F7981: entity F port map(lamdaA => P(7)(981),lamdaB => P(7)(989),lamdaOut => P(6)(981));
U_F7982: entity F port map(lamdaA => P(7)(982),lamdaB => P(7)(990),lamdaOut => P(6)(982));
U_F7983: entity F port map(lamdaA => P(7)(983),lamdaB => P(7)(991),lamdaOut => P(6)(983));
U_G7984: entity G port map(lamdaA => P(7)(976),lamdaB => P(7)(984),s => s(7)(488),lamdaOut => P(6)(984));
U_G7985: entity G port map(lamdaA => P(7)(977),lamdaB => P(7)(985),s => s(7)(489),lamdaOut => P(6)(985));
U_G7986: entity G port map(lamdaA => P(7)(978),lamdaB => P(7)(986),s => s(7)(490),lamdaOut => P(6)(986));
U_G7987: entity G port map(lamdaA => P(7)(979),lamdaB => P(7)(987),s => s(7)(491),lamdaOut => P(6)(987));
U_G7988: entity G port map(lamdaA => P(7)(980),lamdaB => P(7)(988),s => s(7)(492),lamdaOut => P(6)(988));
U_G7989: entity G port map(lamdaA => P(7)(981),lamdaB => P(7)(989),s => s(7)(493),lamdaOut => P(6)(989));
U_G7990: entity G port map(lamdaA => P(7)(982),lamdaB => P(7)(990),s => s(7)(494),lamdaOut => P(6)(990));
U_G7991: entity G port map(lamdaA => P(7)(983),lamdaB => P(7)(991),s => s(7)(495),lamdaOut => P(6)(991));
U_F7992: entity F port map(lamdaA => P(7)(992),lamdaB => P(7)(1000),lamdaOut => P(6)(992));
U_F7993: entity F port map(lamdaA => P(7)(993),lamdaB => P(7)(1001),lamdaOut => P(6)(993));
U_F7994: entity F port map(lamdaA => P(7)(994),lamdaB => P(7)(1002),lamdaOut => P(6)(994));
U_F7995: entity F port map(lamdaA => P(7)(995),lamdaB => P(7)(1003),lamdaOut => P(6)(995));
U_F7996: entity F port map(lamdaA => P(7)(996),lamdaB => P(7)(1004),lamdaOut => P(6)(996));
U_F7997: entity F port map(lamdaA => P(7)(997),lamdaB => P(7)(1005),lamdaOut => P(6)(997));
U_F7998: entity F port map(lamdaA => P(7)(998),lamdaB => P(7)(1006),lamdaOut => P(6)(998));
U_F7999: entity F port map(lamdaA => P(7)(999),lamdaB => P(7)(1007),lamdaOut => P(6)(999));
U_G71000: entity G port map(lamdaA => P(7)(992),lamdaB => P(7)(1000),s => s(7)(496),lamdaOut => P(6)(1000));
U_G71001: entity G port map(lamdaA => P(7)(993),lamdaB => P(7)(1001),s => s(7)(497),lamdaOut => P(6)(1001));
U_G71002: entity G port map(lamdaA => P(7)(994),lamdaB => P(7)(1002),s => s(7)(498),lamdaOut => P(6)(1002));
U_G71003: entity G port map(lamdaA => P(7)(995),lamdaB => P(7)(1003),s => s(7)(499),lamdaOut => P(6)(1003));
U_G71004: entity G port map(lamdaA => P(7)(996),lamdaB => P(7)(1004),s => s(7)(500),lamdaOut => P(6)(1004));
U_G71005: entity G port map(lamdaA => P(7)(997),lamdaB => P(7)(1005),s => s(7)(501),lamdaOut => P(6)(1005));
U_G71006: entity G port map(lamdaA => P(7)(998),lamdaB => P(7)(1006),s => s(7)(502),lamdaOut => P(6)(1006));
U_G71007: entity G port map(lamdaA => P(7)(999),lamdaB => P(7)(1007),s => s(7)(503),lamdaOut => P(6)(1007));
U_F71008: entity F port map(lamdaA => P(7)(1008),lamdaB => P(7)(1016),lamdaOut => P(6)(1008));
U_F71009: entity F port map(lamdaA => P(7)(1009),lamdaB => P(7)(1017),lamdaOut => P(6)(1009));
U_F71010: entity F port map(lamdaA => P(7)(1010),lamdaB => P(7)(1018),lamdaOut => P(6)(1010));
U_F71011: entity F port map(lamdaA => P(7)(1011),lamdaB => P(7)(1019),lamdaOut => P(6)(1011));
U_F71012: entity F port map(lamdaA => P(7)(1012),lamdaB => P(7)(1020),lamdaOut => P(6)(1012));
U_F71013: entity F port map(lamdaA => P(7)(1013),lamdaB => P(7)(1021),lamdaOut => P(6)(1013));
U_F71014: entity F port map(lamdaA => P(7)(1014),lamdaB => P(7)(1022),lamdaOut => P(6)(1014));
U_F71015: entity F port map(lamdaA => P(7)(1015),lamdaB => P(7)(1023),lamdaOut => P(6)(1015));
U_G71016: entity G port map(lamdaA => P(7)(1008),lamdaB => P(7)(1016),s => s(7)(504),lamdaOut => P(6)(1016));
U_G71017: entity G port map(lamdaA => P(7)(1009),lamdaB => P(7)(1017),s => s(7)(505),lamdaOut => P(6)(1017));
U_G71018: entity G port map(lamdaA => P(7)(1010),lamdaB => P(7)(1018),s => s(7)(506),lamdaOut => P(6)(1018));
U_G71019: entity G port map(lamdaA => P(7)(1011),lamdaB => P(7)(1019),s => s(7)(507),lamdaOut => P(6)(1019));
U_G71020: entity G port map(lamdaA => P(7)(1012),lamdaB => P(7)(1020),s => s(7)(508),lamdaOut => P(6)(1020));
U_G71021: entity G port map(lamdaA => P(7)(1013),lamdaB => P(7)(1021),s => s(7)(509),lamdaOut => P(6)(1021));
U_G71022: entity G port map(lamdaA => P(7)(1014),lamdaB => P(7)(1022),s => s(7)(510),lamdaOut => P(6)(1022));
U_G71023: entity G port map(lamdaA => P(7)(1015),lamdaB => P(7)(1023),s => s(7)(511),lamdaOut => P(6)(1023));
-- STAGE 5
U_F60: entity F port map(lamdaA => P(6)(0),lamdaB => P(6)(16),lamdaOut => P(5)(0));
U_F61: entity F port map(lamdaA => P(6)(1),lamdaB => P(6)(17),lamdaOut => P(5)(1));
U_F62: entity F port map(lamdaA => P(6)(2),lamdaB => P(6)(18),lamdaOut => P(5)(2));
U_F63: entity F port map(lamdaA => P(6)(3),lamdaB => P(6)(19),lamdaOut => P(5)(3));
U_F64: entity F port map(lamdaA => P(6)(4),lamdaB => P(6)(20),lamdaOut => P(5)(4));
U_F65: entity F port map(lamdaA => P(6)(5),lamdaB => P(6)(21),lamdaOut => P(5)(5));
U_F66: entity F port map(lamdaA => P(6)(6),lamdaB => P(6)(22),lamdaOut => P(5)(6));
U_F67: entity F port map(lamdaA => P(6)(7),lamdaB => P(6)(23),lamdaOut => P(5)(7));
U_F68: entity F port map(lamdaA => P(6)(8),lamdaB => P(6)(24),lamdaOut => P(5)(8));
U_F69: entity F port map(lamdaA => P(6)(9),lamdaB => P(6)(25),lamdaOut => P(5)(9));
U_F610: entity F port map(lamdaA => P(6)(10),lamdaB => P(6)(26),lamdaOut => P(5)(10));
U_F611: entity F port map(lamdaA => P(6)(11),lamdaB => P(6)(27),lamdaOut => P(5)(11));
U_F612: entity F port map(lamdaA => P(6)(12),lamdaB => P(6)(28),lamdaOut => P(5)(12));
U_F613: entity F port map(lamdaA => P(6)(13),lamdaB => P(6)(29),lamdaOut => P(5)(13));
U_F614: entity F port map(lamdaA => P(6)(14),lamdaB => P(6)(30),lamdaOut => P(5)(14));
U_F615: entity F port map(lamdaA => P(6)(15),lamdaB => P(6)(31),lamdaOut => P(5)(15));
U_G616: entity G port map(lamdaA => P(6)(0),lamdaB => P(6)(16),s => s(6)(0),lamdaOut => P(5)(16));
U_G617: entity G port map(lamdaA => P(6)(1),lamdaB => P(6)(17),s => s(6)(1),lamdaOut => P(5)(17));
U_G618: entity G port map(lamdaA => P(6)(2),lamdaB => P(6)(18),s => s(6)(2),lamdaOut => P(5)(18));
U_G619: entity G port map(lamdaA => P(6)(3),lamdaB => P(6)(19),s => s(6)(3),lamdaOut => P(5)(19));
U_G620: entity G port map(lamdaA => P(6)(4),lamdaB => P(6)(20),s => s(6)(4),lamdaOut => P(5)(20));
U_G621: entity G port map(lamdaA => P(6)(5),lamdaB => P(6)(21),s => s(6)(5),lamdaOut => P(5)(21));
U_G622: entity G port map(lamdaA => P(6)(6),lamdaB => P(6)(22),s => s(6)(6),lamdaOut => P(5)(22));
U_G623: entity G port map(lamdaA => P(6)(7),lamdaB => P(6)(23),s => s(6)(7),lamdaOut => P(5)(23));
U_G624: entity G port map(lamdaA => P(6)(8),lamdaB => P(6)(24),s => s(6)(8),lamdaOut => P(5)(24));
U_G625: entity G port map(lamdaA => P(6)(9),lamdaB => P(6)(25),s => s(6)(9),lamdaOut => P(5)(25));
U_G626: entity G port map(lamdaA => P(6)(10),lamdaB => P(6)(26),s => s(6)(10),lamdaOut => P(5)(26));
U_G627: entity G port map(lamdaA => P(6)(11),lamdaB => P(6)(27),s => s(6)(11),lamdaOut => P(5)(27));
U_G628: entity G port map(lamdaA => P(6)(12),lamdaB => P(6)(28),s => s(6)(12),lamdaOut => P(5)(28));
U_G629: entity G port map(lamdaA => P(6)(13),lamdaB => P(6)(29),s => s(6)(13),lamdaOut => P(5)(29));
U_G630: entity G port map(lamdaA => P(6)(14),lamdaB => P(6)(30),s => s(6)(14),lamdaOut => P(5)(30));
U_G631: entity G port map(lamdaA => P(6)(15),lamdaB => P(6)(31),s => s(6)(15),lamdaOut => P(5)(31));
U_F632: entity F port map(lamdaA => P(6)(32),lamdaB => P(6)(48),lamdaOut => P(5)(32));
U_F633: entity F port map(lamdaA => P(6)(33),lamdaB => P(6)(49),lamdaOut => P(5)(33));
U_F634: entity F port map(lamdaA => P(6)(34),lamdaB => P(6)(50),lamdaOut => P(5)(34));
U_F635: entity F port map(lamdaA => P(6)(35),lamdaB => P(6)(51),lamdaOut => P(5)(35));
U_F636: entity F port map(lamdaA => P(6)(36),lamdaB => P(6)(52),lamdaOut => P(5)(36));
U_F637: entity F port map(lamdaA => P(6)(37),lamdaB => P(6)(53),lamdaOut => P(5)(37));
U_F638: entity F port map(lamdaA => P(6)(38),lamdaB => P(6)(54),lamdaOut => P(5)(38));
U_F639: entity F port map(lamdaA => P(6)(39),lamdaB => P(6)(55),lamdaOut => P(5)(39));
U_F640: entity F port map(lamdaA => P(6)(40),lamdaB => P(6)(56),lamdaOut => P(5)(40));
U_F641: entity F port map(lamdaA => P(6)(41),lamdaB => P(6)(57),lamdaOut => P(5)(41));
U_F642: entity F port map(lamdaA => P(6)(42),lamdaB => P(6)(58),lamdaOut => P(5)(42));
U_F643: entity F port map(lamdaA => P(6)(43),lamdaB => P(6)(59),lamdaOut => P(5)(43));
U_F644: entity F port map(lamdaA => P(6)(44),lamdaB => P(6)(60),lamdaOut => P(5)(44));
U_F645: entity F port map(lamdaA => P(6)(45),lamdaB => P(6)(61),lamdaOut => P(5)(45));
U_F646: entity F port map(lamdaA => P(6)(46),lamdaB => P(6)(62),lamdaOut => P(5)(46));
U_F647: entity F port map(lamdaA => P(6)(47),lamdaB => P(6)(63),lamdaOut => P(5)(47));
U_G648: entity G port map(lamdaA => P(6)(32),lamdaB => P(6)(48),s => s(6)(16),lamdaOut => P(5)(48));
U_G649: entity G port map(lamdaA => P(6)(33),lamdaB => P(6)(49),s => s(6)(17),lamdaOut => P(5)(49));
U_G650: entity G port map(lamdaA => P(6)(34),lamdaB => P(6)(50),s => s(6)(18),lamdaOut => P(5)(50));
U_G651: entity G port map(lamdaA => P(6)(35),lamdaB => P(6)(51),s => s(6)(19),lamdaOut => P(5)(51));
U_G652: entity G port map(lamdaA => P(6)(36),lamdaB => P(6)(52),s => s(6)(20),lamdaOut => P(5)(52));
U_G653: entity G port map(lamdaA => P(6)(37),lamdaB => P(6)(53),s => s(6)(21),lamdaOut => P(5)(53));
U_G654: entity G port map(lamdaA => P(6)(38),lamdaB => P(6)(54),s => s(6)(22),lamdaOut => P(5)(54));
U_G655: entity G port map(lamdaA => P(6)(39),lamdaB => P(6)(55),s => s(6)(23),lamdaOut => P(5)(55));
U_G656: entity G port map(lamdaA => P(6)(40),lamdaB => P(6)(56),s => s(6)(24),lamdaOut => P(5)(56));
U_G657: entity G port map(lamdaA => P(6)(41),lamdaB => P(6)(57),s => s(6)(25),lamdaOut => P(5)(57));
U_G658: entity G port map(lamdaA => P(6)(42),lamdaB => P(6)(58),s => s(6)(26),lamdaOut => P(5)(58));
U_G659: entity G port map(lamdaA => P(6)(43),lamdaB => P(6)(59),s => s(6)(27),lamdaOut => P(5)(59));
U_G660: entity G port map(lamdaA => P(6)(44),lamdaB => P(6)(60),s => s(6)(28),lamdaOut => P(5)(60));
U_G661: entity G port map(lamdaA => P(6)(45),lamdaB => P(6)(61),s => s(6)(29),lamdaOut => P(5)(61));
U_G662: entity G port map(lamdaA => P(6)(46),lamdaB => P(6)(62),s => s(6)(30),lamdaOut => P(5)(62));
U_G663: entity G port map(lamdaA => P(6)(47),lamdaB => P(6)(63),s => s(6)(31),lamdaOut => P(5)(63));
U_F664: entity F port map(lamdaA => P(6)(64),lamdaB => P(6)(80),lamdaOut => P(5)(64));
U_F665: entity F port map(lamdaA => P(6)(65),lamdaB => P(6)(81),lamdaOut => P(5)(65));
U_F666: entity F port map(lamdaA => P(6)(66),lamdaB => P(6)(82),lamdaOut => P(5)(66));
U_F667: entity F port map(lamdaA => P(6)(67),lamdaB => P(6)(83),lamdaOut => P(5)(67));
U_F668: entity F port map(lamdaA => P(6)(68),lamdaB => P(6)(84),lamdaOut => P(5)(68));
U_F669: entity F port map(lamdaA => P(6)(69),lamdaB => P(6)(85),lamdaOut => P(5)(69));
U_F670: entity F port map(lamdaA => P(6)(70),lamdaB => P(6)(86),lamdaOut => P(5)(70));
U_F671: entity F port map(lamdaA => P(6)(71),lamdaB => P(6)(87),lamdaOut => P(5)(71));
U_F672: entity F port map(lamdaA => P(6)(72),lamdaB => P(6)(88),lamdaOut => P(5)(72));
U_F673: entity F port map(lamdaA => P(6)(73),lamdaB => P(6)(89),lamdaOut => P(5)(73));
U_F674: entity F port map(lamdaA => P(6)(74),lamdaB => P(6)(90),lamdaOut => P(5)(74));
U_F675: entity F port map(lamdaA => P(6)(75),lamdaB => P(6)(91),lamdaOut => P(5)(75));
U_F676: entity F port map(lamdaA => P(6)(76),lamdaB => P(6)(92),lamdaOut => P(5)(76));
U_F677: entity F port map(lamdaA => P(6)(77),lamdaB => P(6)(93),lamdaOut => P(5)(77));
U_F678: entity F port map(lamdaA => P(6)(78),lamdaB => P(6)(94),lamdaOut => P(5)(78));
U_F679: entity F port map(lamdaA => P(6)(79),lamdaB => P(6)(95),lamdaOut => P(5)(79));
U_G680: entity G port map(lamdaA => P(6)(64),lamdaB => P(6)(80),s => s(6)(32),lamdaOut => P(5)(80));
U_G681: entity G port map(lamdaA => P(6)(65),lamdaB => P(6)(81),s => s(6)(33),lamdaOut => P(5)(81));
U_G682: entity G port map(lamdaA => P(6)(66),lamdaB => P(6)(82),s => s(6)(34),lamdaOut => P(5)(82));
U_G683: entity G port map(lamdaA => P(6)(67),lamdaB => P(6)(83),s => s(6)(35),lamdaOut => P(5)(83));
U_G684: entity G port map(lamdaA => P(6)(68),lamdaB => P(6)(84),s => s(6)(36),lamdaOut => P(5)(84));
U_G685: entity G port map(lamdaA => P(6)(69),lamdaB => P(6)(85),s => s(6)(37),lamdaOut => P(5)(85));
U_G686: entity G port map(lamdaA => P(6)(70),lamdaB => P(6)(86),s => s(6)(38),lamdaOut => P(5)(86));
U_G687: entity G port map(lamdaA => P(6)(71),lamdaB => P(6)(87),s => s(6)(39),lamdaOut => P(5)(87));
U_G688: entity G port map(lamdaA => P(6)(72),lamdaB => P(6)(88),s => s(6)(40),lamdaOut => P(5)(88));
U_G689: entity G port map(lamdaA => P(6)(73),lamdaB => P(6)(89),s => s(6)(41),lamdaOut => P(5)(89));
U_G690: entity G port map(lamdaA => P(6)(74),lamdaB => P(6)(90),s => s(6)(42),lamdaOut => P(5)(90));
U_G691: entity G port map(lamdaA => P(6)(75),lamdaB => P(6)(91),s => s(6)(43),lamdaOut => P(5)(91));
U_G692: entity G port map(lamdaA => P(6)(76),lamdaB => P(6)(92),s => s(6)(44),lamdaOut => P(5)(92));
U_G693: entity G port map(lamdaA => P(6)(77),lamdaB => P(6)(93),s => s(6)(45),lamdaOut => P(5)(93));
U_G694: entity G port map(lamdaA => P(6)(78),lamdaB => P(6)(94),s => s(6)(46),lamdaOut => P(5)(94));
U_G695: entity G port map(lamdaA => P(6)(79),lamdaB => P(6)(95),s => s(6)(47),lamdaOut => P(5)(95));
U_F696: entity F port map(lamdaA => P(6)(96),lamdaB => P(6)(112),lamdaOut => P(5)(96));
U_F697: entity F port map(lamdaA => P(6)(97),lamdaB => P(6)(113),lamdaOut => P(5)(97));
U_F698: entity F port map(lamdaA => P(6)(98),lamdaB => P(6)(114),lamdaOut => P(5)(98));
U_F699: entity F port map(lamdaA => P(6)(99),lamdaB => P(6)(115),lamdaOut => P(5)(99));
U_F6100: entity F port map(lamdaA => P(6)(100),lamdaB => P(6)(116),lamdaOut => P(5)(100));
U_F6101: entity F port map(lamdaA => P(6)(101),lamdaB => P(6)(117),lamdaOut => P(5)(101));
U_F6102: entity F port map(lamdaA => P(6)(102),lamdaB => P(6)(118),lamdaOut => P(5)(102));
U_F6103: entity F port map(lamdaA => P(6)(103),lamdaB => P(6)(119),lamdaOut => P(5)(103));
U_F6104: entity F port map(lamdaA => P(6)(104),lamdaB => P(6)(120),lamdaOut => P(5)(104));
U_F6105: entity F port map(lamdaA => P(6)(105),lamdaB => P(6)(121),lamdaOut => P(5)(105));
U_F6106: entity F port map(lamdaA => P(6)(106),lamdaB => P(6)(122),lamdaOut => P(5)(106));
U_F6107: entity F port map(lamdaA => P(6)(107),lamdaB => P(6)(123),lamdaOut => P(5)(107));
U_F6108: entity F port map(lamdaA => P(6)(108),lamdaB => P(6)(124),lamdaOut => P(5)(108));
U_F6109: entity F port map(lamdaA => P(6)(109),lamdaB => P(6)(125),lamdaOut => P(5)(109));
U_F6110: entity F port map(lamdaA => P(6)(110),lamdaB => P(6)(126),lamdaOut => P(5)(110));
U_F6111: entity F port map(lamdaA => P(6)(111),lamdaB => P(6)(127),lamdaOut => P(5)(111));
U_G6112: entity G port map(lamdaA => P(6)(96),lamdaB => P(6)(112),s => s(6)(48),lamdaOut => P(5)(112));
U_G6113: entity G port map(lamdaA => P(6)(97),lamdaB => P(6)(113),s => s(6)(49),lamdaOut => P(5)(113));
U_G6114: entity G port map(lamdaA => P(6)(98),lamdaB => P(6)(114),s => s(6)(50),lamdaOut => P(5)(114));
U_G6115: entity G port map(lamdaA => P(6)(99),lamdaB => P(6)(115),s => s(6)(51),lamdaOut => P(5)(115));
U_G6116: entity G port map(lamdaA => P(6)(100),lamdaB => P(6)(116),s => s(6)(52),lamdaOut => P(5)(116));
U_G6117: entity G port map(lamdaA => P(6)(101),lamdaB => P(6)(117),s => s(6)(53),lamdaOut => P(5)(117));
U_G6118: entity G port map(lamdaA => P(6)(102),lamdaB => P(6)(118),s => s(6)(54),lamdaOut => P(5)(118));
U_G6119: entity G port map(lamdaA => P(6)(103),lamdaB => P(6)(119),s => s(6)(55),lamdaOut => P(5)(119));
U_G6120: entity G port map(lamdaA => P(6)(104),lamdaB => P(6)(120),s => s(6)(56),lamdaOut => P(5)(120));
U_G6121: entity G port map(lamdaA => P(6)(105),lamdaB => P(6)(121),s => s(6)(57),lamdaOut => P(5)(121));
U_G6122: entity G port map(lamdaA => P(6)(106),lamdaB => P(6)(122),s => s(6)(58),lamdaOut => P(5)(122));
U_G6123: entity G port map(lamdaA => P(6)(107),lamdaB => P(6)(123),s => s(6)(59),lamdaOut => P(5)(123));
U_G6124: entity G port map(lamdaA => P(6)(108),lamdaB => P(6)(124),s => s(6)(60),lamdaOut => P(5)(124));
U_G6125: entity G port map(lamdaA => P(6)(109),lamdaB => P(6)(125),s => s(6)(61),lamdaOut => P(5)(125));
U_G6126: entity G port map(lamdaA => P(6)(110),lamdaB => P(6)(126),s => s(6)(62),lamdaOut => P(5)(126));
U_G6127: entity G port map(lamdaA => P(6)(111),lamdaB => P(6)(127),s => s(6)(63),lamdaOut => P(5)(127));
U_F6128: entity F port map(lamdaA => P(6)(128),lamdaB => P(6)(144),lamdaOut => P(5)(128));
U_F6129: entity F port map(lamdaA => P(6)(129),lamdaB => P(6)(145),lamdaOut => P(5)(129));
U_F6130: entity F port map(lamdaA => P(6)(130),lamdaB => P(6)(146),lamdaOut => P(5)(130));
U_F6131: entity F port map(lamdaA => P(6)(131),lamdaB => P(6)(147),lamdaOut => P(5)(131));
U_F6132: entity F port map(lamdaA => P(6)(132),lamdaB => P(6)(148),lamdaOut => P(5)(132));
U_F6133: entity F port map(lamdaA => P(6)(133),lamdaB => P(6)(149),lamdaOut => P(5)(133));
U_F6134: entity F port map(lamdaA => P(6)(134),lamdaB => P(6)(150),lamdaOut => P(5)(134));
U_F6135: entity F port map(lamdaA => P(6)(135),lamdaB => P(6)(151),lamdaOut => P(5)(135));
U_F6136: entity F port map(lamdaA => P(6)(136),lamdaB => P(6)(152),lamdaOut => P(5)(136));
U_F6137: entity F port map(lamdaA => P(6)(137),lamdaB => P(6)(153),lamdaOut => P(5)(137));
U_F6138: entity F port map(lamdaA => P(6)(138),lamdaB => P(6)(154),lamdaOut => P(5)(138));
U_F6139: entity F port map(lamdaA => P(6)(139),lamdaB => P(6)(155),lamdaOut => P(5)(139));
U_F6140: entity F port map(lamdaA => P(6)(140),lamdaB => P(6)(156),lamdaOut => P(5)(140));
U_F6141: entity F port map(lamdaA => P(6)(141),lamdaB => P(6)(157),lamdaOut => P(5)(141));
U_F6142: entity F port map(lamdaA => P(6)(142),lamdaB => P(6)(158),lamdaOut => P(5)(142));
U_F6143: entity F port map(lamdaA => P(6)(143),lamdaB => P(6)(159),lamdaOut => P(5)(143));
U_G6144: entity G port map(lamdaA => P(6)(128),lamdaB => P(6)(144),s => s(6)(64),lamdaOut => P(5)(144));
U_G6145: entity G port map(lamdaA => P(6)(129),lamdaB => P(6)(145),s => s(6)(65),lamdaOut => P(5)(145));
U_G6146: entity G port map(lamdaA => P(6)(130),lamdaB => P(6)(146),s => s(6)(66),lamdaOut => P(5)(146));
U_G6147: entity G port map(lamdaA => P(6)(131),lamdaB => P(6)(147),s => s(6)(67),lamdaOut => P(5)(147));
U_G6148: entity G port map(lamdaA => P(6)(132),lamdaB => P(6)(148),s => s(6)(68),lamdaOut => P(5)(148));
U_G6149: entity G port map(lamdaA => P(6)(133),lamdaB => P(6)(149),s => s(6)(69),lamdaOut => P(5)(149));
U_G6150: entity G port map(lamdaA => P(6)(134),lamdaB => P(6)(150),s => s(6)(70),lamdaOut => P(5)(150));
U_G6151: entity G port map(lamdaA => P(6)(135),lamdaB => P(6)(151),s => s(6)(71),lamdaOut => P(5)(151));
U_G6152: entity G port map(lamdaA => P(6)(136),lamdaB => P(6)(152),s => s(6)(72),lamdaOut => P(5)(152));
U_G6153: entity G port map(lamdaA => P(6)(137),lamdaB => P(6)(153),s => s(6)(73),lamdaOut => P(5)(153));
U_G6154: entity G port map(lamdaA => P(6)(138),lamdaB => P(6)(154),s => s(6)(74),lamdaOut => P(5)(154));
U_G6155: entity G port map(lamdaA => P(6)(139),lamdaB => P(6)(155),s => s(6)(75),lamdaOut => P(5)(155));
U_G6156: entity G port map(lamdaA => P(6)(140),lamdaB => P(6)(156),s => s(6)(76),lamdaOut => P(5)(156));
U_G6157: entity G port map(lamdaA => P(6)(141),lamdaB => P(6)(157),s => s(6)(77),lamdaOut => P(5)(157));
U_G6158: entity G port map(lamdaA => P(6)(142),lamdaB => P(6)(158),s => s(6)(78),lamdaOut => P(5)(158));
U_G6159: entity G port map(lamdaA => P(6)(143),lamdaB => P(6)(159),s => s(6)(79),lamdaOut => P(5)(159));
U_F6160: entity F port map(lamdaA => P(6)(160),lamdaB => P(6)(176),lamdaOut => P(5)(160));
U_F6161: entity F port map(lamdaA => P(6)(161),lamdaB => P(6)(177),lamdaOut => P(5)(161));
U_F6162: entity F port map(lamdaA => P(6)(162),lamdaB => P(6)(178),lamdaOut => P(5)(162));
U_F6163: entity F port map(lamdaA => P(6)(163),lamdaB => P(6)(179),lamdaOut => P(5)(163));
U_F6164: entity F port map(lamdaA => P(6)(164),lamdaB => P(6)(180),lamdaOut => P(5)(164));
U_F6165: entity F port map(lamdaA => P(6)(165),lamdaB => P(6)(181),lamdaOut => P(5)(165));
U_F6166: entity F port map(lamdaA => P(6)(166),lamdaB => P(6)(182),lamdaOut => P(5)(166));
U_F6167: entity F port map(lamdaA => P(6)(167),lamdaB => P(6)(183),lamdaOut => P(5)(167));
U_F6168: entity F port map(lamdaA => P(6)(168),lamdaB => P(6)(184),lamdaOut => P(5)(168));
U_F6169: entity F port map(lamdaA => P(6)(169),lamdaB => P(6)(185),lamdaOut => P(5)(169));
U_F6170: entity F port map(lamdaA => P(6)(170),lamdaB => P(6)(186),lamdaOut => P(5)(170));
U_F6171: entity F port map(lamdaA => P(6)(171),lamdaB => P(6)(187),lamdaOut => P(5)(171));
U_F6172: entity F port map(lamdaA => P(6)(172),lamdaB => P(6)(188),lamdaOut => P(5)(172));
U_F6173: entity F port map(lamdaA => P(6)(173),lamdaB => P(6)(189),lamdaOut => P(5)(173));
U_F6174: entity F port map(lamdaA => P(6)(174),lamdaB => P(6)(190),lamdaOut => P(5)(174));
U_F6175: entity F port map(lamdaA => P(6)(175),lamdaB => P(6)(191),lamdaOut => P(5)(175));
U_G6176: entity G port map(lamdaA => P(6)(160),lamdaB => P(6)(176),s => s(6)(80),lamdaOut => P(5)(176));
U_G6177: entity G port map(lamdaA => P(6)(161),lamdaB => P(6)(177),s => s(6)(81),lamdaOut => P(5)(177));
U_G6178: entity G port map(lamdaA => P(6)(162),lamdaB => P(6)(178),s => s(6)(82),lamdaOut => P(5)(178));
U_G6179: entity G port map(lamdaA => P(6)(163),lamdaB => P(6)(179),s => s(6)(83),lamdaOut => P(5)(179));
U_G6180: entity G port map(lamdaA => P(6)(164),lamdaB => P(6)(180),s => s(6)(84),lamdaOut => P(5)(180));
U_G6181: entity G port map(lamdaA => P(6)(165),lamdaB => P(6)(181),s => s(6)(85),lamdaOut => P(5)(181));
U_G6182: entity G port map(lamdaA => P(6)(166),lamdaB => P(6)(182),s => s(6)(86),lamdaOut => P(5)(182));
U_G6183: entity G port map(lamdaA => P(6)(167),lamdaB => P(6)(183),s => s(6)(87),lamdaOut => P(5)(183));
U_G6184: entity G port map(lamdaA => P(6)(168),lamdaB => P(6)(184),s => s(6)(88),lamdaOut => P(5)(184));
U_G6185: entity G port map(lamdaA => P(6)(169),lamdaB => P(6)(185),s => s(6)(89),lamdaOut => P(5)(185));
U_G6186: entity G port map(lamdaA => P(6)(170),lamdaB => P(6)(186),s => s(6)(90),lamdaOut => P(5)(186));
U_G6187: entity G port map(lamdaA => P(6)(171),lamdaB => P(6)(187),s => s(6)(91),lamdaOut => P(5)(187));
U_G6188: entity G port map(lamdaA => P(6)(172),lamdaB => P(6)(188),s => s(6)(92),lamdaOut => P(5)(188));
U_G6189: entity G port map(lamdaA => P(6)(173),lamdaB => P(6)(189),s => s(6)(93),lamdaOut => P(5)(189));
U_G6190: entity G port map(lamdaA => P(6)(174),lamdaB => P(6)(190),s => s(6)(94),lamdaOut => P(5)(190));
U_G6191: entity G port map(lamdaA => P(6)(175),lamdaB => P(6)(191),s => s(6)(95),lamdaOut => P(5)(191));
U_F6192: entity F port map(lamdaA => P(6)(192),lamdaB => P(6)(208),lamdaOut => P(5)(192));
U_F6193: entity F port map(lamdaA => P(6)(193),lamdaB => P(6)(209),lamdaOut => P(5)(193));
U_F6194: entity F port map(lamdaA => P(6)(194),lamdaB => P(6)(210),lamdaOut => P(5)(194));
U_F6195: entity F port map(lamdaA => P(6)(195),lamdaB => P(6)(211),lamdaOut => P(5)(195));
U_F6196: entity F port map(lamdaA => P(6)(196),lamdaB => P(6)(212),lamdaOut => P(5)(196));
U_F6197: entity F port map(lamdaA => P(6)(197),lamdaB => P(6)(213),lamdaOut => P(5)(197));
U_F6198: entity F port map(lamdaA => P(6)(198),lamdaB => P(6)(214),lamdaOut => P(5)(198));
U_F6199: entity F port map(lamdaA => P(6)(199),lamdaB => P(6)(215),lamdaOut => P(5)(199));
U_F6200: entity F port map(lamdaA => P(6)(200),lamdaB => P(6)(216),lamdaOut => P(5)(200));
U_F6201: entity F port map(lamdaA => P(6)(201),lamdaB => P(6)(217),lamdaOut => P(5)(201));
U_F6202: entity F port map(lamdaA => P(6)(202),lamdaB => P(6)(218),lamdaOut => P(5)(202));
U_F6203: entity F port map(lamdaA => P(6)(203),lamdaB => P(6)(219),lamdaOut => P(5)(203));
U_F6204: entity F port map(lamdaA => P(6)(204),lamdaB => P(6)(220),lamdaOut => P(5)(204));
U_F6205: entity F port map(lamdaA => P(6)(205),lamdaB => P(6)(221),lamdaOut => P(5)(205));
U_F6206: entity F port map(lamdaA => P(6)(206),lamdaB => P(6)(222),lamdaOut => P(5)(206));
U_F6207: entity F port map(lamdaA => P(6)(207),lamdaB => P(6)(223),lamdaOut => P(5)(207));
U_G6208: entity G port map(lamdaA => P(6)(192),lamdaB => P(6)(208),s => s(6)(96),lamdaOut => P(5)(208));
U_G6209: entity G port map(lamdaA => P(6)(193),lamdaB => P(6)(209),s => s(6)(97),lamdaOut => P(5)(209));
U_G6210: entity G port map(lamdaA => P(6)(194),lamdaB => P(6)(210),s => s(6)(98),lamdaOut => P(5)(210));
U_G6211: entity G port map(lamdaA => P(6)(195),lamdaB => P(6)(211),s => s(6)(99),lamdaOut => P(5)(211));
U_G6212: entity G port map(lamdaA => P(6)(196),lamdaB => P(6)(212),s => s(6)(100),lamdaOut => P(5)(212));
U_G6213: entity G port map(lamdaA => P(6)(197),lamdaB => P(6)(213),s => s(6)(101),lamdaOut => P(5)(213));
U_G6214: entity G port map(lamdaA => P(6)(198),lamdaB => P(6)(214),s => s(6)(102),lamdaOut => P(5)(214));
U_G6215: entity G port map(lamdaA => P(6)(199),lamdaB => P(6)(215),s => s(6)(103),lamdaOut => P(5)(215));
U_G6216: entity G port map(lamdaA => P(6)(200),lamdaB => P(6)(216),s => s(6)(104),lamdaOut => P(5)(216));
U_G6217: entity G port map(lamdaA => P(6)(201),lamdaB => P(6)(217),s => s(6)(105),lamdaOut => P(5)(217));
U_G6218: entity G port map(lamdaA => P(6)(202),lamdaB => P(6)(218),s => s(6)(106),lamdaOut => P(5)(218));
U_G6219: entity G port map(lamdaA => P(6)(203),lamdaB => P(6)(219),s => s(6)(107),lamdaOut => P(5)(219));
U_G6220: entity G port map(lamdaA => P(6)(204),lamdaB => P(6)(220),s => s(6)(108),lamdaOut => P(5)(220));
U_G6221: entity G port map(lamdaA => P(6)(205),lamdaB => P(6)(221),s => s(6)(109),lamdaOut => P(5)(221));
U_G6222: entity G port map(lamdaA => P(6)(206),lamdaB => P(6)(222),s => s(6)(110),lamdaOut => P(5)(222));
U_G6223: entity G port map(lamdaA => P(6)(207),lamdaB => P(6)(223),s => s(6)(111),lamdaOut => P(5)(223));
U_F6224: entity F port map(lamdaA => P(6)(224),lamdaB => P(6)(240),lamdaOut => P(5)(224));
U_F6225: entity F port map(lamdaA => P(6)(225),lamdaB => P(6)(241),lamdaOut => P(5)(225));
U_F6226: entity F port map(lamdaA => P(6)(226),lamdaB => P(6)(242),lamdaOut => P(5)(226));
U_F6227: entity F port map(lamdaA => P(6)(227),lamdaB => P(6)(243),lamdaOut => P(5)(227));
U_F6228: entity F port map(lamdaA => P(6)(228),lamdaB => P(6)(244),lamdaOut => P(5)(228));
U_F6229: entity F port map(lamdaA => P(6)(229),lamdaB => P(6)(245),lamdaOut => P(5)(229));
U_F6230: entity F port map(lamdaA => P(6)(230),lamdaB => P(6)(246),lamdaOut => P(5)(230));
U_F6231: entity F port map(lamdaA => P(6)(231),lamdaB => P(6)(247),lamdaOut => P(5)(231));
U_F6232: entity F port map(lamdaA => P(6)(232),lamdaB => P(6)(248),lamdaOut => P(5)(232));
U_F6233: entity F port map(lamdaA => P(6)(233),lamdaB => P(6)(249),lamdaOut => P(5)(233));
U_F6234: entity F port map(lamdaA => P(6)(234),lamdaB => P(6)(250),lamdaOut => P(5)(234));
U_F6235: entity F port map(lamdaA => P(6)(235),lamdaB => P(6)(251),lamdaOut => P(5)(235));
U_F6236: entity F port map(lamdaA => P(6)(236),lamdaB => P(6)(252),lamdaOut => P(5)(236));
U_F6237: entity F port map(lamdaA => P(6)(237),lamdaB => P(6)(253),lamdaOut => P(5)(237));
U_F6238: entity F port map(lamdaA => P(6)(238),lamdaB => P(6)(254),lamdaOut => P(5)(238));
U_F6239: entity F port map(lamdaA => P(6)(239),lamdaB => P(6)(255),lamdaOut => P(5)(239));
U_G6240: entity G port map(lamdaA => P(6)(224),lamdaB => P(6)(240),s => s(6)(112),lamdaOut => P(5)(240));
U_G6241: entity G port map(lamdaA => P(6)(225),lamdaB => P(6)(241),s => s(6)(113),lamdaOut => P(5)(241));
U_G6242: entity G port map(lamdaA => P(6)(226),lamdaB => P(6)(242),s => s(6)(114),lamdaOut => P(5)(242));
U_G6243: entity G port map(lamdaA => P(6)(227),lamdaB => P(6)(243),s => s(6)(115),lamdaOut => P(5)(243));
U_G6244: entity G port map(lamdaA => P(6)(228),lamdaB => P(6)(244),s => s(6)(116),lamdaOut => P(5)(244));
U_G6245: entity G port map(lamdaA => P(6)(229),lamdaB => P(6)(245),s => s(6)(117),lamdaOut => P(5)(245));
U_G6246: entity G port map(lamdaA => P(6)(230),lamdaB => P(6)(246),s => s(6)(118),lamdaOut => P(5)(246));
U_G6247: entity G port map(lamdaA => P(6)(231),lamdaB => P(6)(247),s => s(6)(119),lamdaOut => P(5)(247));
U_G6248: entity G port map(lamdaA => P(6)(232),lamdaB => P(6)(248),s => s(6)(120),lamdaOut => P(5)(248));
U_G6249: entity G port map(lamdaA => P(6)(233),lamdaB => P(6)(249),s => s(6)(121),lamdaOut => P(5)(249));
U_G6250: entity G port map(lamdaA => P(6)(234),lamdaB => P(6)(250),s => s(6)(122),lamdaOut => P(5)(250));
U_G6251: entity G port map(lamdaA => P(6)(235),lamdaB => P(6)(251),s => s(6)(123),lamdaOut => P(5)(251));
U_G6252: entity G port map(lamdaA => P(6)(236),lamdaB => P(6)(252),s => s(6)(124),lamdaOut => P(5)(252));
U_G6253: entity G port map(lamdaA => P(6)(237),lamdaB => P(6)(253),s => s(6)(125),lamdaOut => P(5)(253));
U_G6254: entity G port map(lamdaA => P(6)(238),lamdaB => P(6)(254),s => s(6)(126),lamdaOut => P(5)(254));
U_G6255: entity G port map(lamdaA => P(6)(239),lamdaB => P(6)(255),s => s(6)(127),lamdaOut => P(5)(255));
U_F6256: entity F port map(lamdaA => P(6)(256),lamdaB => P(6)(272),lamdaOut => P(5)(256));
U_F6257: entity F port map(lamdaA => P(6)(257),lamdaB => P(6)(273),lamdaOut => P(5)(257));
U_F6258: entity F port map(lamdaA => P(6)(258),lamdaB => P(6)(274),lamdaOut => P(5)(258));
U_F6259: entity F port map(lamdaA => P(6)(259),lamdaB => P(6)(275),lamdaOut => P(5)(259));
U_F6260: entity F port map(lamdaA => P(6)(260),lamdaB => P(6)(276),lamdaOut => P(5)(260));
U_F6261: entity F port map(lamdaA => P(6)(261),lamdaB => P(6)(277),lamdaOut => P(5)(261));
U_F6262: entity F port map(lamdaA => P(6)(262),lamdaB => P(6)(278),lamdaOut => P(5)(262));
U_F6263: entity F port map(lamdaA => P(6)(263),lamdaB => P(6)(279),lamdaOut => P(5)(263));
U_F6264: entity F port map(lamdaA => P(6)(264),lamdaB => P(6)(280),lamdaOut => P(5)(264));
U_F6265: entity F port map(lamdaA => P(6)(265),lamdaB => P(6)(281),lamdaOut => P(5)(265));
U_F6266: entity F port map(lamdaA => P(6)(266),lamdaB => P(6)(282),lamdaOut => P(5)(266));
U_F6267: entity F port map(lamdaA => P(6)(267),lamdaB => P(6)(283),lamdaOut => P(5)(267));
U_F6268: entity F port map(lamdaA => P(6)(268),lamdaB => P(6)(284),lamdaOut => P(5)(268));
U_F6269: entity F port map(lamdaA => P(6)(269),lamdaB => P(6)(285),lamdaOut => P(5)(269));
U_F6270: entity F port map(lamdaA => P(6)(270),lamdaB => P(6)(286),lamdaOut => P(5)(270));
U_F6271: entity F port map(lamdaA => P(6)(271),lamdaB => P(6)(287),lamdaOut => P(5)(271));
U_G6272: entity G port map(lamdaA => P(6)(256),lamdaB => P(6)(272),s => s(6)(128),lamdaOut => P(5)(272));
U_G6273: entity G port map(lamdaA => P(6)(257),lamdaB => P(6)(273),s => s(6)(129),lamdaOut => P(5)(273));
U_G6274: entity G port map(lamdaA => P(6)(258),lamdaB => P(6)(274),s => s(6)(130),lamdaOut => P(5)(274));
U_G6275: entity G port map(lamdaA => P(6)(259),lamdaB => P(6)(275),s => s(6)(131),lamdaOut => P(5)(275));
U_G6276: entity G port map(lamdaA => P(6)(260),lamdaB => P(6)(276),s => s(6)(132),lamdaOut => P(5)(276));
U_G6277: entity G port map(lamdaA => P(6)(261),lamdaB => P(6)(277),s => s(6)(133),lamdaOut => P(5)(277));
U_G6278: entity G port map(lamdaA => P(6)(262),lamdaB => P(6)(278),s => s(6)(134),lamdaOut => P(5)(278));
U_G6279: entity G port map(lamdaA => P(6)(263),lamdaB => P(6)(279),s => s(6)(135),lamdaOut => P(5)(279));
U_G6280: entity G port map(lamdaA => P(6)(264),lamdaB => P(6)(280),s => s(6)(136),lamdaOut => P(5)(280));
U_G6281: entity G port map(lamdaA => P(6)(265),lamdaB => P(6)(281),s => s(6)(137),lamdaOut => P(5)(281));
U_G6282: entity G port map(lamdaA => P(6)(266),lamdaB => P(6)(282),s => s(6)(138),lamdaOut => P(5)(282));
U_G6283: entity G port map(lamdaA => P(6)(267),lamdaB => P(6)(283),s => s(6)(139),lamdaOut => P(5)(283));
U_G6284: entity G port map(lamdaA => P(6)(268),lamdaB => P(6)(284),s => s(6)(140),lamdaOut => P(5)(284));
U_G6285: entity G port map(lamdaA => P(6)(269),lamdaB => P(6)(285),s => s(6)(141),lamdaOut => P(5)(285));
U_G6286: entity G port map(lamdaA => P(6)(270),lamdaB => P(6)(286),s => s(6)(142),lamdaOut => P(5)(286));
U_G6287: entity G port map(lamdaA => P(6)(271),lamdaB => P(6)(287),s => s(6)(143),lamdaOut => P(5)(287));
U_F6288: entity F port map(lamdaA => P(6)(288),lamdaB => P(6)(304),lamdaOut => P(5)(288));
U_F6289: entity F port map(lamdaA => P(6)(289),lamdaB => P(6)(305),lamdaOut => P(5)(289));
U_F6290: entity F port map(lamdaA => P(6)(290),lamdaB => P(6)(306),lamdaOut => P(5)(290));
U_F6291: entity F port map(lamdaA => P(6)(291),lamdaB => P(6)(307),lamdaOut => P(5)(291));
U_F6292: entity F port map(lamdaA => P(6)(292),lamdaB => P(6)(308),lamdaOut => P(5)(292));
U_F6293: entity F port map(lamdaA => P(6)(293),lamdaB => P(6)(309),lamdaOut => P(5)(293));
U_F6294: entity F port map(lamdaA => P(6)(294),lamdaB => P(6)(310),lamdaOut => P(5)(294));
U_F6295: entity F port map(lamdaA => P(6)(295),lamdaB => P(6)(311),lamdaOut => P(5)(295));
U_F6296: entity F port map(lamdaA => P(6)(296),lamdaB => P(6)(312),lamdaOut => P(5)(296));
U_F6297: entity F port map(lamdaA => P(6)(297),lamdaB => P(6)(313),lamdaOut => P(5)(297));
U_F6298: entity F port map(lamdaA => P(6)(298),lamdaB => P(6)(314),lamdaOut => P(5)(298));
U_F6299: entity F port map(lamdaA => P(6)(299),lamdaB => P(6)(315),lamdaOut => P(5)(299));
U_F6300: entity F port map(lamdaA => P(6)(300),lamdaB => P(6)(316),lamdaOut => P(5)(300));
U_F6301: entity F port map(lamdaA => P(6)(301),lamdaB => P(6)(317),lamdaOut => P(5)(301));
U_F6302: entity F port map(lamdaA => P(6)(302),lamdaB => P(6)(318),lamdaOut => P(5)(302));
U_F6303: entity F port map(lamdaA => P(6)(303),lamdaB => P(6)(319),lamdaOut => P(5)(303));
U_G6304: entity G port map(lamdaA => P(6)(288),lamdaB => P(6)(304),s => s(6)(144),lamdaOut => P(5)(304));
U_G6305: entity G port map(lamdaA => P(6)(289),lamdaB => P(6)(305),s => s(6)(145),lamdaOut => P(5)(305));
U_G6306: entity G port map(lamdaA => P(6)(290),lamdaB => P(6)(306),s => s(6)(146),lamdaOut => P(5)(306));
U_G6307: entity G port map(lamdaA => P(6)(291),lamdaB => P(6)(307),s => s(6)(147),lamdaOut => P(5)(307));
U_G6308: entity G port map(lamdaA => P(6)(292),lamdaB => P(6)(308),s => s(6)(148),lamdaOut => P(5)(308));
U_G6309: entity G port map(lamdaA => P(6)(293),lamdaB => P(6)(309),s => s(6)(149),lamdaOut => P(5)(309));
U_G6310: entity G port map(lamdaA => P(6)(294),lamdaB => P(6)(310),s => s(6)(150),lamdaOut => P(5)(310));
U_G6311: entity G port map(lamdaA => P(6)(295),lamdaB => P(6)(311),s => s(6)(151),lamdaOut => P(5)(311));
U_G6312: entity G port map(lamdaA => P(6)(296),lamdaB => P(6)(312),s => s(6)(152),lamdaOut => P(5)(312));
U_G6313: entity G port map(lamdaA => P(6)(297),lamdaB => P(6)(313),s => s(6)(153),lamdaOut => P(5)(313));
U_G6314: entity G port map(lamdaA => P(6)(298),lamdaB => P(6)(314),s => s(6)(154),lamdaOut => P(5)(314));
U_G6315: entity G port map(lamdaA => P(6)(299),lamdaB => P(6)(315),s => s(6)(155),lamdaOut => P(5)(315));
U_G6316: entity G port map(lamdaA => P(6)(300),lamdaB => P(6)(316),s => s(6)(156),lamdaOut => P(5)(316));
U_G6317: entity G port map(lamdaA => P(6)(301),lamdaB => P(6)(317),s => s(6)(157),lamdaOut => P(5)(317));
U_G6318: entity G port map(lamdaA => P(6)(302),lamdaB => P(6)(318),s => s(6)(158),lamdaOut => P(5)(318));
U_G6319: entity G port map(lamdaA => P(6)(303),lamdaB => P(6)(319),s => s(6)(159),lamdaOut => P(5)(319));
U_F6320: entity F port map(lamdaA => P(6)(320),lamdaB => P(6)(336),lamdaOut => P(5)(320));
U_F6321: entity F port map(lamdaA => P(6)(321),lamdaB => P(6)(337),lamdaOut => P(5)(321));
U_F6322: entity F port map(lamdaA => P(6)(322),lamdaB => P(6)(338),lamdaOut => P(5)(322));
U_F6323: entity F port map(lamdaA => P(6)(323),lamdaB => P(6)(339),lamdaOut => P(5)(323));
U_F6324: entity F port map(lamdaA => P(6)(324),lamdaB => P(6)(340),lamdaOut => P(5)(324));
U_F6325: entity F port map(lamdaA => P(6)(325),lamdaB => P(6)(341),lamdaOut => P(5)(325));
U_F6326: entity F port map(lamdaA => P(6)(326),lamdaB => P(6)(342),lamdaOut => P(5)(326));
U_F6327: entity F port map(lamdaA => P(6)(327),lamdaB => P(6)(343),lamdaOut => P(5)(327));
U_F6328: entity F port map(lamdaA => P(6)(328),lamdaB => P(6)(344),lamdaOut => P(5)(328));
U_F6329: entity F port map(lamdaA => P(6)(329),lamdaB => P(6)(345),lamdaOut => P(5)(329));
U_F6330: entity F port map(lamdaA => P(6)(330),lamdaB => P(6)(346),lamdaOut => P(5)(330));
U_F6331: entity F port map(lamdaA => P(6)(331),lamdaB => P(6)(347),lamdaOut => P(5)(331));
U_F6332: entity F port map(lamdaA => P(6)(332),lamdaB => P(6)(348),lamdaOut => P(5)(332));
U_F6333: entity F port map(lamdaA => P(6)(333),lamdaB => P(6)(349),lamdaOut => P(5)(333));
U_F6334: entity F port map(lamdaA => P(6)(334),lamdaB => P(6)(350),lamdaOut => P(5)(334));
U_F6335: entity F port map(lamdaA => P(6)(335),lamdaB => P(6)(351),lamdaOut => P(5)(335));
U_G6336: entity G port map(lamdaA => P(6)(320),lamdaB => P(6)(336),s => s(6)(160),lamdaOut => P(5)(336));
U_G6337: entity G port map(lamdaA => P(6)(321),lamdaB => P(6)(337),s => s(6)(161),lamdaOut => P(5)(337));
U_G6338: entity G port map(lamdaA => P(6)(322),lamdaB => P(6)(338),s => s(6)(162),lamdaOut => P(5)(338));
U_G6339: entity G port map(lamdaA => P(6)(323),lamdaB => P(6)(339),s => s(6)(163),lamdaOut => P(5)(339));
U_G6340: entity G port map(lamdaA => P(6)(324),lamdaB => P(6)(340),s => s(6)(164),lamdaOut => P(5)(340));
U_G6341: entity G port map(lamdaA => P(6)(325),lamdaB => P(6)(341),s => s(6)(165),lamdaOut => P(5)(341));
U_G6342: entity G port map(lamdaA => P(6)(326),lamdaB => P(6)(342),s => s(6)(166),lamdaOut => P(5)(342));
U_G6343: entity G port map(lamdaA => P(6)(327),lamdaB => P(6)(343),s => s(6)(167),lamdaOut => P(5)(343));
U_G6344: entity G port map(lamdaA => P(6)(328),lamdaB => P(6)(344),s => s(6)(168),lamdaOut => P(5)(344));
U_G6345: entity G port map(lamdaA => P(6)(329),lamdaB => P(6)(345),s => s(6)(169),lamdaOut => P(5)(345));
U_G6346: entity G port map(lamdaA => P(6)(330),lamdaB => P(6)(346),s => s(6)(170),lamdaOut => P(5)(346));
U_G6347: entity G port map(lamdaA => P(6)(331),lamdaB => P(6)(347),s => s(6)(171),lamdaOut => P(5)(347));
U_G6348: entity G port map(lamdaA => P(6)(332),lamdaB => P(6)(348),s => s(6)(172),lamdaOut => P(5)(348));
U_G6349: entity G port map(lamdaA => P(6)(333),lamdaB => P(6)(349),s => s(6)(173),lamdaOut => P(5)(349));
U_G6350: entity G port map(lamdaA => P(6)(334),lamdaB => P(6)(350),s => s(6)(174),lamdaOut => P(5)(350));
U_G6351: entity G port map(lamdaA => P(6)(335),lamdaB => P(6)(351),s => s(6)(175),lamdaOut => P(5)(351));
U_F6352: entity F port map(lamdaA => P(6)(352),lamdaB => P(6)(368),lamdaOut => P(5)(352));
U_F6353: entity F port map(lamdaA => P(6)(353),lamdaB => P(6)(369),lamdaOut => P(5)(353));
U_F6354: entity F port map(lamdaA => P(6)(354),lamdaB => P(6)(370),lamdaOut => P(5)(354));
U_F6355: entity F port map(lamdaA => P(6)(355),lamdaB => P(6)(371),lamdaOut => P(5)(355));
U_F6356: entity F port map(lamdaA => P(6)(356),lamdaB => P(6)(372),lamdaOut => P(5)(356));
U_F6357: entity F port map(lamdaA => P(6)(357),lamdaB => P(6)(373),lamdaOut => P(5)(357));
U_F6358: entity F port map(lamdaA => P(6)(358),lamdaB => P(6)(374),lamdaOut => P(5)(358));
U_F6359: entity F port map(lamdaA => P(6)(359),lamdaB => P(6)(375),lamdaOut => P(5)(359));
U_F6360: entity F port map(lamdaA => P(6)(360),lamdaB => P(6)(376),lamdaOut => P(5)(360));
U_F6361: entity F port map(lamdaA => P(6)(361),lamdaB => P(6)(377),lamdaOut => P(5)(361));
U_F6362: entity F port map(lamdaA => P(6)(362),lamdaB => P(6)(378),lamdaOut => P(5)(362));
U_F6363: entity F port map(lamdaA => P(6)(363),lamdaB => P(6)(379),lamdaOut => P(5)(363));
U_F6364: entity F port map(lamdaA => P(6)(364),lamdaB => P(6)(380),lamdaOut => P(5)(364));
U_F6365: entity F port map(lamdaA => P(6)(365),lamdaB => P(6)(381),lamdaOut => P(5)(365));
U_F6366: entity F port map(lamdaA => P(6)(366),lamdaB => P(6)(382),lamdaOut => P(5)(366));
U_F6367: entity F port map(lamdaA => P(6)(367),lamdaB => P(6)(383),lamdaOut => P(5)(367));
U_G6368: entity G port map(lamdaA => P(6)(352),lamdaB => P(6)(368),s => s(6)(176),lamdaOut => P(5)(368));
U_G6369: entity G port map(lamdaA => P(6)(353),lamdaB => P(6)(369),s => s(6)(177),lamdaOut => P(5)(369));
U_G6370: entity G port map(lamdaA => P(6)(354),lamdaB => P(6)(370),s => s(6)(178),lamdaOut => P(5)(370));
U_G6371: entity G port map(lamdaA => P(6)(355),lamdaB => P(6)(371),s => s(6)(179),lamdaOut => P(5)(371));
U_G6372: entity G port map(lamdaA => P(6)(356),lamdaB => P(6)(372),s => s(6)(180),lamdaOut => P(5)(372));
U_G6373: entity G port map(lamdaA => P(6)(357),lamdaB => P(6)(373),s => s(6)(181),lamdaOut => P(5)(373));
U_G6374: entity G port map(lamdaA => P(6)(358),lamdaB => P(6)(374),s => s(6)(182),lamdaOut => P(5)(374));
U_G6375: entity G port map(lamdaA => P(6)(359),lamdaB => P(6)(375),s => s(6)(183),lamdaOut => P(5)(375));
U_G6376: entity G port map(lamdaA => P(6)(360),lamdaB => P(6)(376),s => s(6)(184),lamdaOut => P(5)(376));
U_G6377: entity G port map(lamdaA => P(6)(361),lamdaB => P(6)(377),s => s(6)(185),lamdaOut => P(5)(377));
U_G6378: entity G port map(lamdaA => P(6)(362),lamdaB => P(6)(378),s => s(6)(186),lamdaOut => P(5)(378));
U_G6379: entity G port map(lamdaA => P(6)(363),lamdaB => P(6)(379),s => s(6)(187),lamdaOut => P(5)(379));
U_G6380: entity G port map(lamdaA => P(6)(364),lamdaB => P(6)(380),s => s(6)(188),lamdaOut => P(5)(380));
U_G6381: entity G port map(lamdaA => P(6)(365),lamdaB => P(6)(381),s => s(6)(189),lamdaOut => P(5)(381));
U_G6382: entity G port map(lamdaA => P(6)(366),lamdaB => P(6)(382),s => s(6)(190),lamdaOut => P(5)(382));
U_G6383: entity G port map(lamdaA => P(6)(367),lamdaB => P(6)(383),s => s(6)(191),lamdaOut => P(5)(383));
U_F6384: entity F port map(lamdaA => P(6)(384),lamdaB => P(6)(400),lamdaOut => P(5)(384));
U_F6385: entity F port map(lamdaA => P(6)(385),lamdaB => P(6)(401),lamdaOut => P(5)(385));
U_F6386: entity F port map(lamdaA => P(6)(386),lamdaB => P(6)(402),lamdaOut => P(5)(386));
U_F6387: entity F port map(lamdaA => P(6)(387),lamdaB => P(6)(403),lamdaOut => P(5)(387));
U_F6388: entity F port map(lamdaA => P(6)(388),lamdaB => P(6)(404),lamdaOut => P(5)(388));
U_F6389: entity F port map(lamdaA => P(6)(389),lamdaB => P(6)(405),lamdaOut => P(5)(389));
U_F6390: entity F port map(lamdaA => P(6)(390),lamdaB => P(6)(406),lamdaOut => P(5)(390));
U_F6391: entity F port map(lamdaA => P(6)(391),lamdaB => P(6)(407),lamdaOut => P(5)(391));
U_F6392: entity F port map(lamdaA => P(6)(392),lamdaB => P(6)(408),lamdaOut => P(5)(392));
U_F6393: entity F port map(lamdaA => P(6)(393),lamdaB => P(6)(409),lamdaOut => P(5)(393));
U_F6394: entity F port map(lamdaA => P(6)(394),lamdaB => P(6)(410),lamdaOut => P(5)(394));
U_F6395: entity F port map(lamdaA => P(6)(395),lamdaB => P(6)(411),lamdaOut => P(5)(395));
U_F6396: entity F port map(lamdaA => P(6)(396),lamdaB => P(6)(412),lamdaOut => P(5)(396));
U_F6397: entity F port map(lamdaA => P(6)(397),lamdaB => P(6)(413),lamdaOut => P(5)(397));
U_F6398: entity F port map(lamdaA => P(6)(398),lamdaB => P(6)(414),lamdaOut => P(5)(398));
U_F6399: entity F port map(lamdaA => P(6)(399),lamdaB => P(6)(415),lamdaOut => P(5)(399));
U_G6400: entity G port map(lamdaA => P(6)(384),lamdaB => P(6)(400),s => s(6)(192),lamdaOut => P(5)(400));
U_G6401: entity G port map(lamdaA => P(6)(385),lamdaB => P(6)(401),s => s(6)(193),lamdaOut => P(5)(401));
U_G6402: entity G port map(lamdaA => P(6)(386),lamdaB => P(6)(402),s => s(6)(194),lamdaOut => P(5)(402));
U_G6403: entity G port map(lamdaA => P(6)(387),lamdaB => P(6)(403),s => s(6)(195),lamdaOut => P(5)(403));
U_G6404: entity G port map(lamdaA => P(6)(388),lamdaB => P(6)(404),s => s(6)(196),lamdaOut => P(5)(404));
U_G6405: entity G port map(lamdaA => P(6)(389),lamdaB => P(6)(405),s => s(6)(197),lamdaOut => P(5)(405));
U_G6406: entity G port map(lamdaA => P(6)(390),lamdaB => P(6)(406),s => s(6)(198),lamdaOut => P(5)(406));
U_G6407: entity G port map(lamdaA => P(6)(391),lamdaB => P(6)(407),s => s(6)(199),lamdaOut => P(5)(407));
U_G6408: entity G port map(lamdaA => P(6)(392),lamdaB => P(6)(408),s => s(6)(200),lamdaOut => P(5)(408));
U_G6409: entity G port map(lamdaA => P(6)(393),lamdaB => P(6)(409),s => s(6)(201),lamdaOut => P(5)(409));
U_G6410: entity G port map(lamdaA => P(6)(394),lamdaB => P(6)(410),s => s(6)(202),lamdaOut => P(5)(410));
U_G6411: entity G port map(lamdaA => P(6)(395),lamdaB => P(6)(411),s => s(6)(203),lamdaOut => P(5)(411));
U_G6412: entity G port map(lamdaA => P(6)(396),lamdaB => P(6)(412),s => s(6)(204),lamdaOut => P(5)(412));
U_G6413: entity G port map(lamdaA => P(6)(397),lamdaB => P(6)(413),s => s(6)(205),lamdaOut => P(5)(413));
U_G6414: entity G port map(lamdaA => P(6)(398),lamdaB => P(6)(414),s => s(6)(206),lamdaOut => P(5)(414));
U_G6415: entity G port map(lamdaA => P(6)(399),lamdaB => P(6)(415),s => s(6)(207),lamdaOut => P(5)(415));
U_F6416: entity F port map(lamdaA => P(6)(416),lamdaB => P(6)(432),lamdaOut => P(5)(416));
U_F6417: entity F port map(lamdaA => P(6)(417),lamdaB => P(6)(433),lamdaOut => P(5)(417));
U_F6418: entity F port map(lamdaA => P(6)(418),lamdaB => P(6)(434),lamdaOut => P(5)(418));
U_F6419: entity F port map(lamdaA => P(6)(419),lamdaB => P(6)(435),lamdaOut => P(5)(419));
U_F6420: entity F port map(lamdaA => P(6)(420),lamdaB => P(6)(436),lamdaOut => P(5)(420));
U_F6421: entity F port map(lamdaA => P(6)(421),lamdaB => P(6)(437),lamdaOut => P(5)(421));
U_F6422: entity F port map(lamdaA => P(6)(422),lamdaB => P(6)(438),lamdaOut => P(5)(422));
U_F6423: entity F port map(lamdaA => P(6)(423),lamdaB => P(6)(439),lamdaOut => P(5)(423));
U_F6424: entity F port map(lamdaA => P(6)(424),lamdaB => P(6)(440),lamdaOut => P(5)(424));
U_F6425: entity F port map(lamdaA => P(6)(425),lamdaB => P(6)(441),lamdaOut => P(5)(425));
U_F6426: entity F port map(lamdaA => P(6)(426),lamdaB => P(6)(442),lamdaOut => P(5)(426));
U_F6427: entity F port map(lamdaA => P(6)(427),lamdaB => P(6)(443),lamdaOut => P(5)(427));
U_F6428: entity F port map(lamdaA => P(6)(428),lamdaB => P(6)(444),lamdaOut => P(5)(428));
U_F6429: entity F port map(lamdaA => P(6)(429),lamdaB => P(6)(445),lamdaOut => P(5)(429));
U_F6430: entity F port map(lamdaA => P(6)(430),lamdaB => P(6)(446),lamdaOut => P(5)(430));
U_F6431: entity F port map(lamdaA => P(6)(431),lamdaB => P(6)(447),lamdaOut => P(5)(431));
U_G6432: entity G port map(lamdaA => P(6)(416),lamdaB => P(6)(432),s => s(6)(208),lamdaOut => P(5)(432));
U_G6433: entity G port map(lamdaA => P(6)(417),lamdaB => P(6)(433),s => s(6)(209),lamdaOut => P(5)(433));
U_G6434: entity G port map(lamdaA => P(6)(418),lamdaB => P(6)(434),s => s(6)(210),lamdaOut => P(5)(434));
U_G6435: entity G port map(lamdaA => P(6)(419),lamdaB => P(6)(435),s => s(6)(211),lamdaOut => P(5)(435));
U_G6436: entity G port map(lamdaA => P(6)(420),lamdaB => P(6)(436),s => s(6)(212),lamdaOut => P(5)(436));
U_G6437: entity G port map(lamdaA => P(6)(421),lamdaB => P(6)(437),s => s(6)(213),lamdaOut => P(5)(437));
U_G6438: entity G port map(lamdaA => P(6)(422),lamdaB => P(6)(438),s => s(6)(214),lamdaOut => P(5)(438));
U_G6439: entity G port map(lamdaA => P(6)(423),lamdaB => P(6)(439),s => s(6)(215),lamdaOut => P(5)(439));
U_G6440: entity G port map(lamdaA => P(6)(424),lamdaB => P(6)(440),s => s(6)(216),lamdaOut => P(5)(440));
U_G6441: entity G port map(lamdaA => P(6)(425),lamdaB => P(6)(441),s => s(6)(217),lamdaOut => P(5)(441));
U_G6442: entity G port map(lamdaA => P(6)(426),lamdaB => P(6)(442),s => s(6)(218),lamdaOut => P(5)(442));
U_G6443: entity G port map(lamdaA => P(6)(427),lamdaB => P(6)(443),s => s(6)(219),lamdaOut => P(5)(443));
U_G6444: entity G port map(lamdaA => P(6)(428),lamdaB => P(6)(444),s => s(6)(220),lamdaOut => P(5)(444));
U_G6445: entity G port map(lamdaA => P(6)(429),lamdaB => P(6)(445),s => s(6)(221),lamdaOut => P(5)(445));
U_G6446: entity G port map(lamdaA => P(6)(430),lamdaB => P(6)(446),s => s(6)(222),lamdaOut => P(5)(446));
U_G6447: entity G port map(lamdaA => P(6)(431),lamdaB => P(6)(447),s => s(6)(223),lamdaOut => P(5)(447));
U_F6448: entity F port map(lamdaA => P(6)(448),lamdaB => P(6)(464),lamdaOut => P(5)(448));
U_F6449: entity F port map(lamdaA => P(6)(449),lamdaB => P(6)(465),lamdaOut => P(5)(449));
U_F6450: entity F port map(lamdaA => P(6)(450),lamdaB => P(6)(466),lamdaOut => P(5)(450));
U_F6451: entity F port map(lamdaA => P(6)(451),lamdaB => P(6)(467),lamdaOut => P(5)(451));
U_F6452: entity F port map(lamdaA => P(6)(452),lamdaB => P(6)(468),lamdaOut => P(5)(452));
U_F6453: entity F port map(lamdaA => P(6)(453),lamdaB => P(6)(469),lamdaOut => P(5)(453));
U_F6454: entity F port map(lamdaA => P(6)(454),lamdaB => P(6)(470),lamdaOut => P(5)(454));
U_F6455: entity F port map(lamdaA => P(6)(455),lamdaB => P(6)(471),lamdaOut => P(5)(455));
U_F6456: entity F port map(lamdaA => P(6)(456),lamdaB => P(6)(472),lamdaOut => P(5)(456));
U_F6457: entity F port map(lamdaA => P(6)(457),lamdaB => P(6)(473),lamdaOut => P(5)(457));
U_F6458: entity F port map(lamdaA => P(6)(458),lamdaB => P(6)(474),lamdaOut => P(5)(458));
U_F6459: entity F port map(lamdaA => P(6)(459),lamdaB => P(6)(475),lamdaOut => P(5)(459));
U_F6460: entity F port map(lamdaA => P(6)(460),lamdaB => P(6)(476),lamdaOut => P(5)(460));
U_F6461: entity F port map(lamdaA => P(6)(461),lamdaB => P(6)(477),lamdaOut => P(5)(461));
U_F6462: entity F port map(lamdaA => P(6)(462),lamdaB => P(6)(478),lamdaOut => P(5)(462));
U_F6463: entity F port map(lamdaA => P(6)(463),lamdaB => P(6)(479),lamdaOut => P(5)(463));
U_G6464: entity G port map(lamdaA => P(6)(448),lamdaB => P(6)(464),s => s(6)(224),lamdaOut => P(5)(464));
U_G6465: entity G port map(lamdaA => P(6)(449),lamdaB => P(6)(465),s => s(6)(225),lamdaOut => P(5)(465));
U_G6466: entity G port map(lamdaA => P(6)(450),lamdaB => P(6)(466),s => s(6)(226),lamdaOut => P(5)(466));
U_G6467: entity G port map(lamdaA => P(6)(451),lamdaB => P(6)(467),s => s(6)(227),lamdaOut => P(5)(467));
U_G6468: entity G port map(lamdaA => P(6)(452),lamdaB => P(6)(468),s => s(6)(228),lamdaOut => P(5)(468));
U_G6469: entity G port map(lamdaA => P(6)(453),lamdaB => P(6)(469),s => s(6)(229),lamdaOut => P(5)(469));
U_G6470: entity G port map(lamdaA => P(6)(454),lamdaB => P(6)(470),s => s(6)(230),lamdaOut => P(5)(470));
U_G6471: entity G port map(lamdaA => P(6)(455),lamdaB => P(6)(471),s => s(6)(231),lamdaOut => P(5)(471));
U_G6472: entity G port map(lamdaA => P(6)(456),lamdaB => P(6)(472),s => s(6)(232),lamdaOut => P(5)(472));
U_G6473: entity G port map(lamdaA => P(6)(457),lamdaB => P(6)(473),s => s(6)(233),lamdaOut => P(5)(473));
U_G6474: entity G port map(lamdaA => P(6)(458),lamdaB => P(6)(474),s => s(6)(234),lamdaOut => P(5)(474));
U_G6475: entity G port map(lamdaA => P(6)(459),lamdaB => P(6)(475),s => s(6)(235),lamdaOut => P(5)(475));
U_G6476: entity G port map(lamdaA => P(6)(460),lamdaB => P(6)(476),s => s(6)(236),lamdaOut => P(5)(476));
U_G6477: entity G port map(lamdaA => P(6)(461),lamdaB => P(6)(477),s => s(6)(237),lamdaOut => P(5)(477));
U_G6478: entity G port map(lamdaA => P(6)(462),lamdaB => P(6)(478),s => s(6)(238),lamdaOut => P(5)(478));
U_G6479: entity G port map(lamdaA => P(6)(463),lamdaB => P(6)(479),s => s(6)(239),lamdaOut => P(5)(479));
U_F6480: entity F port map(lamdaA => P(6)(480),lamdaB => P(6)(496),lamdaOut => P(5)(480));
U_F6481: entity F port map(lamdaA => P(6)(481),lamdaB => P(6)(497),lamdaOut => P(5)(481));
U_F6482: entity F port map(lamdaA => P(6)(482),lamdaB => P(6)(498),lamdaOut => P(5)(482));
U_F6483: entity F port map(lamdaA => P(6)(483),lamdaB => P(6)(499),lamdaOut => P(5)(483));
U_F6484: entity F port map(lamdaA => P(6)(484),lamdaB => P(6)(500),lamdaOut => P(5)(484));
U_F6485: entity F port map(lamdaA => P(6)(485),lamdaB => P(6)(501),lamdaOut => P(5)(485));
U_F6486: entity F port map(lamdaA => P(6)(486),lamdaB => P(6)(502),lamdaOut => P(5)(486));
U_F6487: entity F port map(lamdaA => P(6)(487),lamdaB => P(6)(503),lamdaOut => P(5)(487));
U_F6488: entity F port map(lamdaA => P(6)(488),lamdaB => P(6)(504),lamdaOut => P(5)(488));
U_F6489: entity F port map(lamdaA => P(6)(489),lamdaB => P(6)(505),lamdaOut => P(5)(489));
U_F6490: entity F port map(lamdaA => P(6)(490),lamdaB => P(6)(506),lamdaOut => P(5)(490));
U_F6491: entity F port map(lamdaA => P(6)(491),lamdaB => P(6)(507),lamdaOut => P(5)(491));
U_F6492: entity F port map(lamdaA => P(6)(492),lamdaB => P(6)(508),lamdaOut => P(5)(492));
U_F6493: entity F port map(lamdaA => P(6)(493),lamdaB => P(6)(509),lamdaOut => P(5)(493));
U_F6494: entity F port map(lamdaA => P(6)(494),lamdaB => P(6)(510),lamdaOut => P(5)(494));
U_F6495: entity F port map(lamdaA => P(6)(495),lamdaB => P(6)(511),lamdaOut => P(5)(495));
U_G6496: entity G port map(lamdaA => P(6)(480),lamdaB => P(6)(496),s => s(6)(240),lamdaOut => P(5)(496));
U_G6497: entity G port map(lamdaA => P(6)(481),lamdaB => P(6)(497),s => s(6)(241),lamdaOut => P(5)(497));
U_G6498: entity G port map(lamdaA => P(6)(482),lamdaB => P(6)(498),s => s(6)(242),lamdaOut => P(5)(498));
U_G6499: entity G port map(lamdaA => P(6)(483),lamdaB => P(6)(499),s => s(6)(243),lamdaOut => P(5)(499));
U_G6500: entity G port map(lamdaA => P(6)(484),lamdaB => P(6)(500),s => s(6)(244),lamdaOut => P(5)(500));
U_G6501: entity G port map(lamdaA => P(6)(485),lamdaB => P(6)(501),s => s(6)(245),lamdaOut => P(5)(501));
U_G6502: entity G port map(lamdaA => P(6)(486),lamdaB => P(6)(502),s => s(6)(246),lamdaOut => P(5)(502));
U_G6503: entity G port map(lamdaA => P(6)(487),lamdaB => P(6)(503),s => s(6)(247),lamdaOut => P(5)(503));
U_G6504: entity G port map(lamdaA => P(6)(488),lamdaB => P(6)(504),s => s(6)(248),lamdaOut => P(5)(504));
U_G6505: entity G port map(lamdaA => P(6)(489),lamdaB => P(6)(505),s => s(6)(249),lamdaOut => P(5)(505));
U_G6506: entity G port map(lamdaA => P(6)(490),lamdaB => P(6)(506),s => s(6)(250),lamdaOut => P(5)(506));
U_G6507: entity G port map(lamdaA => P(6)(491),lamdaB => P(6)(507),s => s(6)(251),lamdaOut => P(5)(507));
U_G6508: entity G port map(lamdaA => P(6)(492),lamdaB => P(6)(508),s => s(6)(252),lamdaOut => P(5)(508));
U_G6509: entity G port map(lamdaA => P(6)(493),lamdaB => P(6)(509),s => s(6)(253),lamdaOut => P(5)(509));
U_G6510: entity G port map(lamdaA => P(6)(494),lamdaB => P(6)(510),s => s(6)(254),lamdaOut => P(5)(510));
U_G6511: entity G port map(lamdaA => P(6)(495),lamdaB => P(6)(511),s => s(6)(255),lamdaOut => P(5)(511));
U_F6512: entity F port map(lamdaA => P(6)(512),lamdaB => P(6)(528),lamdaOut => P(5)(512));
U_F6513: entity F port map(lamdaA => P(6)(513),lamdaB => P(6)(529),lamdaOut => P(5)(513));
U_F6514: entity F port map(lamdaA => P(6)(514),lamdaB => P(6)(530),lamdaOut => P(5)(514));
U_F6515: entity F port map(lamdaA => P(6)(515),lamdaB => P(6)(531),lamdaOut => P(5)(515));
U_F6516: entity F port map(lamdaA => P(6)(516),lamdaB => P(6)(532),lamdaOut => P(5)(516));
U_F6517: entity F port map(lamdaA => P(6)(517),lamdaB => P(6)(533),lamdaOut => P(5)(517));
U_F6518: entity F port map(lamdaA => P(6)(518),lamdaB => P(6)(534),lamdaOut => P(5)(518));
U_F6519: entity F port map(lamdaA => P(6)(519),lamdaB => P(6)(535),lamdaOut => P(5)(519));
U_F6520: entity F port map(lamdaA => P(6)(520),lamdaB => P(6)(536),lamdaOut => P(5)(520));
U_F6521: entity F port map(lamdaA => P(6)(521),lamdaB => P(6)(537),lamdaOut => P(5)(521));
U_F6522: entity F port map(lamdaA => P(6)(522),lamdaB => P(6)(538),lamdaOut => P(5)(522));
U_F6523: entity F port map(lamdaA => P(6)(523),lamdaB => P(6)(539),lamdaOut => P(5)(523));
U_F6524: entity F port map(lamdaA => P(6)(524),lamdaB => P(6)(540),lamdaOut => P(5)(524));
U_F6525: entity F port map(lamdaA => P(6)(525),lamdaB => P(6)(541),lamdaOut => P(5)(525));
U_F6526: entity F port map(lamdaA => P(6)(526),lamdaB => P(6)(542),lamdaOut => P(5)(526));
U_F6527: entity F port map(lamdaA => P(6)(527),lamdaB => P(6)(543),lamdaOut => P(5)(527));
U_G6528: entity G port map(lamdaA => P(6)(512),lamdaB => P(6)(528),s => s(6)(256),lamdaOut => P(5)(528));
U_G6529: entity G port map(lamdaA => P(6)(513),lamdaB => P(6)(529),s => s(6)(257),lamdaOut => P(5)(529));
U_G6530: entity G port map(lamdaA => P(6)(514),lamdaB => P(6)(530),s => s(6)(258),lamdaOut => P(5)(530));
U_G6531: entity G port map(lamdaA => P(6)(515),lamdaB => P(6)(531),s => s(6)(259),lamdaOut => P(5)(531));
U_G6532: entity G port map(lamdaA => P(6)(516),lamdaB => P(6)(532),s => s(6)(260),lamdaOut => P(5)(532));
U_G6533: entity G port map(lamdaA => P(6)(517),lamdaB => P(6)(533),s => s(6)(261),lamdaOut => P(5)(533));
U_G6534: entity G port map(lamdaA => P(6)(518),lamdaB => P(6)(534),s => s(6)(262),lamdaOut => P(5)(534));
U_G6535: entity G port map(lamdaA => P(6)(519),lamdaB => P(6)(535),s => s(6)(263),lamdaOut => P(5)(535));
U_G6536: entity G port map(lamdaA => P(6)(520),lamdaB => P(6)(536),s => s(6)(264),lamdaOut => P(5)(536));
U_G6537: entity G port map(lamdaA => P(6)(521),lamdaB => P(6)(537),s => s(6)(265),lamdaOut => P(5)(537));
U_G6538: entity G port map(lamdaA => P(6)(522),lamdaB => P(6)(538),s => s(6)(266),lamdaOut => P(5)(538));
U_G6539: entity G port map(lamdaA => P(6)(523),lamdaB => P(6)(539),s => s(6)(267),lamdaOut => P(5)(539));
U_G6540: entity G port map(lamdaA => P(6)(524),lamdaB => P(6)(540),s => s(6)(268),lamdaOut => P(5)(540));
U_G6541: entity G port map(lamdaA => P(6)(525),lamdaB => P(6)(541),s => s(6)(269),lamdaOut => P(5)(541));
U_G6542: entity G port map(lamdaA => P(6)(526),lamdaB => P(6)(542),s => s(6)(270),lamdaOut => P(5)(542));
U_G6543: entity G port map(lamdaA => P(6)(527),lamdaB => P(6)(543),s => s(6)(271),lamdaOut => P(5)(543));
U_F6544: entity F port map(lamdaA => P(6)(544),lamdaB => P(6)(560),lamdaOut => P(5)(544));
U_F6545: entity F port map(lamdaA => P(6)(545),lamdaB => P(6)(561),lamdaOut => P(5)(545));
U_F6546: entity F port map(lamdaA => P(6)(546),lamdaB => P(6)(562),lamdaOut => P(5)(546));
U_F6547: entity F port map(lamdaA => P(6)(547),lamdaB => P(6)(563),lamdaOut => P(5)(547));
U_F6548: entity F port map(lamdaA => P(6)(548),lamdaB => P(6)(564),lamdaOut => P(5)(548));
U_F6549: entity F port map(lamdaA => P(6)(549),lamdaB => P(6)(565),lamdaOut => P(5)(549));
U_F6550: entity F port map(lamdaA => P(6)(550),lamdaB => P(6)(566),lamdaOut => P(5)(550));
U_F6551: entity F port map(lamdaA => P(6)(551),lamdaB => P(6)(567),lamdaOut => P(5)(551));
U_F6552: entity F port map(lamdaA => P(6)(552),lamdaB => P(6)(568),lamdaOut => P(5)(552));
U_F6553: entity F port map(lamdaA => P(6)(553),lamdaB => P(6)(569),lamdaOut => P(5)(553));
U_F6554: entity F port map(lamdaA => P(6)(554),lamdaB => P(6)(570),lamdaOut => P(5)(554));
U_F6555: entity F port map(lamdaA => P(6)(555),lamdaB => P(6)(571),lamdaOut => P(5)(555));
U_F6556: entity F port map(lamdaA => P(6)(556),lamdaB => P(6)(572),lamdaOut => P(5)(556));
U_F6557: entity F port map(lamdaA => P(6)(557),lamdaB => P(6)(573),lamdaOut => P(5)(557));
U_F6558: entity F port map(lamdaA => P(6)(558),lamdaB => P(6)(574),lamdaOut => P(5)(558));
U_F6559: entity F port map(lamdaA => P(6)(559),lamdaB => P(6)(575),lamdaOut => P(5)(559));
U_G6560: entity G port map(lamdaA => P(6)(544),lamdaB => P(6)(560),s => s(6)(272),lamdaOut => P(5)(560));
U_G6561: entity G port map(lamdaA => P(6)(545),lamdaB => P(6)(561),s => s(6)(273),lamdaOut => P(5)(561));
U_G6562: entity G port map(lamdaA => P(6)(546),lamdaB => P(6)(562),s => s(6)(274),lamdaOut => P(5)(562));
U_G6563: entity G port map(lamdaA => P(6)(547),lamdaB => P(6)(563),s => s(6)(275),lamdaOut => P(5)(563));
U_G6564: entity G port map(lamdaA => P(6)(548),lamdaB => P(6)(564),s => s(6)(276),lamdaOut => P(5)(564));
U_G6565: entity G port map(lamdaA => P(6)(549),lamdaB => P(6)(565),s => s(6)(277),lamdaOut => P(5)(565));
U_G6566: entity G port map(lamdaA => P(6)(550),lamdaB => P(6)(566),s => s(6)(278),lamdaOut => P(5)(566));
U_G6567: entity G port map(lamdaA => P(6)(551),lamdaB => P(6)(567),s => s(6)(279),lamdaOut => P(5)(567));
U_G6568: entity G port map(lamdaA => P(6)(552),lamdaB => P(6)(568),s => s(6)(280),lamdaOut => P(5)(568));
U_G6569: entity G port map(lamdaA => P(6)(553),lamdaB => P(6)(569),s => s(6)(281),lamdaOut => P(5)(569));
U_G6570: entity G port map(lamdaA => P(6)(554),lamdaB => P(6)(570),s => s(6)(282),lamdaOut => P(5)(570));
U_G6571: entity G port map(lamdaA => P(6)(555),lamdaB => P(6)(571),s => s(6)(283),lamdaOut => P(5)(571));
U_G6572: entity G port map(lamdaA => P(6)(556),lamdaB => P(6)(572),s => s(6)(284),lamdaOut => P(5)(572));
U_G6573: entity G port map(lamdaA => P(6)(557),lamdaB => P(6)(573),s => s(6)(285),lamdaOut => P(5)(573));
U_G6574: entity G port map(lamdaA => P(6)(558),lamdaB => P(6)(574),s => s(6)(286),lamdaOut => P(5)(574));
U_G6575: entity G port map(lamdaA => P(6)(559),lamdaB => P(6)(575),s => s(6)(287),lamdaOut => P(5)(575));
U_F6576: entity F port map(lamdaA => P(6)(576),lamdaB => P(6)(592),lamdaOut => P(5)(576));
U_F6577: entity F port map(lamdaA => P(6)(577),lamdaB => P(6)(593),lamdaOut => P(5)(577));
U_F6578: entity F port map(lamdaA => P(6)(578),lamdaB => P(6)(594),lamdaOut => P(5)(578));
U_F6579: entity F port map(lamdaA => P(6)(579),lamdaB => P(6)(595),lamdaOut => P(5)(579));
U_F6580: entity F port map(lamdaA => P(6)(580),lamdaB => P(6)(596),lamdaOut => P(5)(580));
U_F6581: entity F port map(lamdaA => P(6)(581),lamdaB => P(6)(597),lamdaOut => P(5)(581));
U_F6582: entity F port map(lamdaA => P(6)(582),lamdaB => P(6)(598),lamdaOut => P(5)(582));
U_F6583: entity F port map(lamdaA => P(6)(583),lamdaB => P(6)(599),lamdaOut => P(5)(583));
U_F6584: entity F port map(lamdaA => P(6)(584),lamdaB => P(6)(600),lamdaOut => P(5)(584));
U_F6585: entity F port map(lamdaA => P(6)(585),lamdaB => P(6)(601),lamdaOut => P(5)(585));
U_F6586: entity F port map(lamdaA => P(6)(586),lamdaB => P(6)(602),lamdaOut => P(5)(586));
U_F6587: entity F port map(lamdaA => P(6)(587),lamdaB => P(6)(603),lamdaOut => P(5)(587));
U_F6588: entity F port map(lamdaA => P(6)(588),lamdaB => P(6)(604),lamdaOut => P(5)(588));
U_F6589: entity F port map(lamdaA => P(6)(589),lamdaB => P(6)(605),lamdaOut => P(5)(589));
U_F6590: entity F port map(lamdaA => P(6)(590),lamdaB => P(6)(606),lamdaOut => P(5)(590));
U_F6591: entity F port map(lamdaA => P(6)(591),lamdaB => P(6)(607),lamdaOut => P(5)(591));
U_G6592: entity G port map(lamdaA => P(6)(576),lamdaB => P(6)(592),s => s(6)(288),lamdaOut => P(5)(592));
U_G6593: entity G port map(lamdaA => P(6)(577),lamdaB => P(6)(593),s => s(6)(289),lamdaOut => P(5)(593));
U_G6594: entity G port map(lamdaA => P(6)(578),lamdaB => P(6)(594),s => s(6)(290),lamdaOut => P(5)(594));
U_G6595: entity G port map(lamdaA => P(6)(579),lamdaB => P(6)(595),s => s(6)(291),lamdaOut => P(5)(595));
U_G6596: entity G port map(lamdaA => P(6)(580),lamdaB => P(6)(596),s => s(6)(292),lamdaOut => P(5)(596));
U_G6597: entity G port map(lamdaA => P(6)(581),lamdaB => P(6)(597),s => s(6)(293),lamdaOut => P(5)(597));
U_G6598: entity G port map(lamdaA => P(6)(582),lamdaB => P(6)(598),s => s(6)(294),lamdaOut => P(5)(598));
U_G6599: entity G port map(lamdaA => P(6)(583),lamdaB => P(6)(599),s => s(6)(295),lamdaOut => P(5)(599));
U_G6600: entity G port map(lamdaA => P(6)(584),lamdaB => P(6)(600),s => s(6)(296),lamdaOut => P(5)(600));
U_G6601: entity G port map(lamdaA => P(6)(585),lamdaB => P(6)(601),s => s(6)(297),lamdaOut => P(5)(601));
U_G6602: entity G port map(lamdaA => P(6)(586),lamdaB => P(6)(602),s => s(6)(298),lamdaOut => P(5)(602));
U_G6603: entity G port map(lamdaA => P(6)(587),lamdaB => P(6)(603),s => s(6)(299),lamdaOut => P(5)(603));
U_G6604: entity G port map(lamdaA => P(6)(588),lamdaB => P(6)(604),s => s(6)(300),lamdaOut => P(5)(604));
U_G6605: entity G port map(lamdaA => P(6)(589),lamdaB => P(6)(605),s => s(6)(301),lamdaOut => P(5)(605));
U_G6606: entity G port map(lamdaA => P(6)(590),lamdaB => P(6)(606),s => s(6)(302),lamdaOut => P(5)(606));
U_G6607: entity G port map(lamdaA => P(6)(591),lamdaB => P(6)(607),s => s(6)(303),lamdaOut => P(5)(607));
U_F6608: entity F port map(lamdaA => P(6)(608),lamdaB => P(6)(624),lamdaOut => P(5)(608));
U_F6609: entity F port map(lamdaA => P(6)(609),lamdaB => P(6)(625),lamdaOut => P(5)(609));
U_F6610: entity F port map(lamdaA => P(6)(610),lamdaB => P(6)(626),lamdaOut => P(5)(610));
U_F6611: entity F port map(lamdaA => P(6)(611),lamdaB => P(6)(627),lamdaOut => P(5)(611));
U_F6612: entity F port map(lamdaA => P(6)(612),lamdaB => P(6)(628),lamdaOut => P(5)(612));
U_F6613: entity F port map(lamdaA => P(6)(613),lamdaB => P(6)(629),lamdaOut => P(5)(613));
U_F6614: entity F port map(lamdaA => P(6)(614),lamdaB => P(6)(630),lamdaOut => P(5)(614));
U_F6615: entity F port map(lamdaA => P(6)(615),lamdaB => P(6)(631),lamdaOut => P(5)(615));
U_F6616: entity F port map(lamdaA => P(6)(616),lamdaB => P(6)(632),lamdaOut => P(5)(616));
U_F6617: entity F port map(lamdaA => P(6)(617),lamdaB => P(6)(633),lamdaOut => P(5)(617));
U_F6618: entity F port map(lamdaA => P(6)(618),lamdaB => P(6)(634),lamdaOut => P(5)(618));
U_F6619: entity F port map(lamdaA => P(6)(619),lamdaB => P(6)(635),lamdaOut => P(5)(619));
U_F6620: entity F port map(lamdaA => P(6)(620),lamdaB => P(6)(636),lamdaOut => P(5)(620));
U_F6621: entity F port map(lamdaA => P(6)(621),lamdaB => P(6)(637),lamdaOut => P(5)(621));
U_F6622: entity F port map(lamdaA => P(6)(622),lamdaB => P(6)(638),lamdaOut => P(5)(622));
U_F6623: entity F port map(lamdaA => P(6)(623),lamdaB => P(6)(639),lamdaOut => P(5)(623));
U_G6624: entity G port map(lamdaA => P(6)(608),lamdaB => P(6)(624),s => s(6)(304),lamdaOut => P(5)(624));
U_G6625: entity G port map(lamdaA => P(6)(609),lamdaB => P(6)(625),s => s(6)(305),lamdaOut => P(5)(625));
U_G6626: entity G port map(lamdaA => P(6)(610),lamdaB => P(6)(626),s => s(6)(306),lamdaOut => P(5)(626));
U_G6627: entity G port map(lamdaA => P(6)(611),lamdaB => P(6)(627),s => s(6)(307),lamdaOut => P(5)(627));
U_G6628: entity G port map(lamdaA => P(6)(612),lamdaB => P(6)(628),s => s(6)(308),lamdaOut => P(5)(628));
U_G6629: entity G port map(lamdaA => P(6)(613),lamdaB => P(6)(629),s => s(6)(309),lamdaOut => P(5)(629));
U_G6630: entity G port map(lamdaA => P(6)(614),lamdaB => P(6)(630),s => s(6)(310),lamdaOut => P(5)(630));
U_G6631: entity G port map(lamdaA => P(6)(615),lamdaB => P(6)(631),s => s(6)(311),lamdaOut => P(5)(631));
U_G6632: entity G port map(lamdaA => P(6)(616),lamdaB => P(6)(632),s => s(6)(312),lamdaOut => P(5)(632));
U_G6633: entity G port map(lamdaA => P(6)(617),lamdaB => P(6)(633),s => s(6)(313),lamdaOut => P(5)(633));
U_G6634: entity G port map(lamdaA => P(6)(618),lamdaB => P(6)(634),s => s(6)(314),lamdaOut => P(5)(634));
U_G6635: entity G port map(lamdaA => P(6)(619),lamdaB => P(6)(635),s => s(6)(315),lamdaOut => P(5)(635));
U_G6636: entity G port map(lamdaA => P(6)(620),lamdaB => P(6)(636),s => s(6)(316),lamdaOut => P(5)(636));
U_G6637: entity G port map(lamdaA => P(6)(621),lamdaB => P(6)(637),s => s(6)(317),lamdaOut => P(5)(637));
U_G6638: entity G port map(lamdaA => P(6)(622),lamdaB => P(6)(638),s => s(6)(318),lamdaOut => P(5)(638));
U_G6639: entity G port map(lamdaA => P(6)(623),lamdaB => P(6)(639),s => s(6)(319),lamdaOut => P(5)(639));
U_F6640: entity F port map(lamdaA => P(6)(640),lamdaB => P(6)(656),lamdaOut => P(5)(640));
U_F6641: entity F port map(lamdaA => P(6)(641),lamdaB => P(6)(657),lamdaOut => P(5)(641));
U_F6642: entity F port map(lamdaA => P(6)(642),lamdaB => P(6)(658),lamdaOut => P(5)(642));
U_F6643: entity F port map(lamdaA => P(6)(643),lamdaB => P(6)(659),lamdaOut => P(5)(643));
U_F6644: entity F port map(lamdaA => P(6)(644),lamdaB => P(6)(660),lamdaOut => P(5)(644));
U_F6645: entity F port map(lamdaA => P(6)(645),lamdaB => P(6)(661),lamdaOut => P(5)(645));
U_F6646: entity F port map(lamdaA => P(6)(646),lamdaB => P(6)(662),lamdaOut => P(5)(646));
U_F6647: entity F port map(lamdaA => P(6)(647),lamdaB => P(6)(663),lamdaOut => P(5)(647));
U_F6648: entity F port map(lamdaA => P(6)(648),lamdaB => P(6)(664),lamdaOut => P(5)(648));
U_F6649: entity F port map(lamdaA => P(6)(649),lamdaB => P(6)(665),lamdaOut => P(5)(649));
U_F6650: entity F port map(lamdaA => P(6)(650),lamdaB => P(6)(666),lamdaOut => P(5)(650));
U_F6651: entity F port map(lamdaA => P(6)(651),lamdaB => P(6)(667),lamdaOut => P(5)(651));
U_F6652: entity F port map(lamdaA => P(6)(652),lamdaB => P(6)(668),lamdaOut => P(5)(652));
U_F6653: entity F port map(lamdaA => P(6)(653),lamdaB => P(6)(669),lamdaOut => P(5)(653));
U_F6654: entity F port map(lamdaA => P(6)(654),lamdaB => P(6)(670),lamdaOut => P(5)(654));
U_F6655: entity F port map(lamdaA => P(6)(655),lamdaB => P(6)(671),lamdaOut => P(5)(655));
U_G6656: entity G port map(lamdaA => P(6)(640),lamdaB => P(6)(656),s => s(6)(320),lamdaOut => P(5)(656));
U_G6657: entity G port map(lamdaA => P(6)(641),lamdaB => P(6)(657),s => s(6)(321),lamdaOut => P(5)(657));
U_G6658: entity G port map(lamdaA => P(6)(642),lamdaB => P(6)(658),s => s(6)(322),lamdaOut => P(5)(658));
U_G6659: entity G port map(lamdaA => P(6)(643),lamdaB => P(6)(659),s => s(6)(323),lamdaOut => P(5)(659));
U_G6660: entity G port map(lamdaA => P(6)(644),lamdaB => P(6)(660),s => s(6)(324),lamdaOut => P(5)(660));
U_G6661: entity G port map(lamdaA => P(6)(645),lamdaB => P(6)(661),s => s(6)(325),lamdaOut => P(5)(661));
U_G6662: entity G port map(lamdaA => P(6)(646),lamdaB => P(6)(662),s => s(6)(326),lamdaOut => P(5)(662));
U_G6663: entity G port map(lamdaA => P(6)(647),lamdaB => P(6)(663),s => s(6)(327),lamdaOut => P(5)(663));
U_G6664: entity G port map(lamdaA => P(6)(648),lamdaB => P(6)(664),s => s(6)(328),lamdaOut => P(5)(664));
U_G6665: entity G port map(lamdaA => P(6)(649),lamdaB => P(6)(665),s => s(6)(329),lamdaOut => P(5)(665));
U_G6666: entity G port map(lamdaA => P(6)(650),lamdaB => P(6)(666),s => s(6)(330),lamdaOut => P(5)(666));
U_G6667: entity G port map(lamdaA => P(6)(651),lamdaB => P(6)(667),s => s(6)(331),lamdaOut => P(5)(667));
U_G6668: entity G port map(lamdaA => P(6)(652),lamdaB => P(6)(668),s => s(6)(332),lamdaOut => P(5)(668));
U_G6669: entity G port map(lamdaA => P(6)(653),lamdaB => P(6)(669),s => s(6)(333),lamdaOut => P(5)(669));
U_G6670: entity G port map(lamdaA => P(6)(654),lamdaB => P(6)(670),s => s(6)(334),lamdaOut => P(5)(670));
U_G6671: entity G port map(lamdaA => P(6)(655),lamdaB => P(6)(671),s => s(6)(335),lamdaOut => P(5)(671));
U_F6672: entity F port map(lamdaA => P(6)(672),lamdaB => P(6)(688),lamdaOut => P(5)(672));
U_F6673: entity F port map(lamdaA => P(6)(673),lamdaB => P(6)(689),lamdaOut => P(5)(673));
U_F6674: entity F port map(lamdaA => P(6)(674),lamdaB => P(6)(690),lamdaOut => P(5)(674));
U_F6675: entity F port map(lamdaA => P(6)(675),lamdaB => P(6)(691),lamdaOut => P(5)(675));
U_F6676: entity F port map(lamdaA => P(6)(676),lamdaB => P(6)(692),lamdaOut => P(5)(676));
U_F6677: entity F port map(lamdaA => P(6)(677),lamdaB => P(6)(693),lamdaOut => P(5)(677));
U_F6678: entity F port map(lamdaA => P(6)(678),lamdaB => P(6)(694),lamdaOut => P(5)(678));
U_F6679: entity F port map(lamdaA => P(6)(679),lamdaB => P(6)(695),lamdaOut => P(5)(679));
U_F6680: entity F port map(lamdaA => P(6)(680),lamdaB => P(6)(696),lamdaOut => P(5)(680));
U_F6681: entity F port map(lamdaA => P(6)(681),lamdaB => P(6)(697),lamdaOut => P(5)(681));
U_F6682: entity F port map(lamdaA => P(6)(682),lamdaB => P(6)(698),lamdaOut => P(5)(682));
U_F6683: entity F port map(lamdaA => P(6)(683),lamdaB => P(6)(699),lamdaOut => P(5)(683));
U_F6684: entity F port map(lamdaA => P(6)(684),lamdaB => P(6)(700),lamdaOut => P(5)(684));
U_F6685: entity F port map(lamdaA => P(6)(685),lamdaB => P(6)(701),lamdaOut => P(5)(685));
U_F6686: entity F port map(lamdaA => P(6)(686),lamdaB => P(6)(702),lamdaOut => P(5)(686));
U_F6687: entity F port map(lamdaA => P(6)(687),lamdaB => P(6)(703),lamdaOut => P(5)(687));
U_G6688: entity G port map(lamdaA => P(6)(672),lamdaB => P(6)(688),s => s(6)(336),lamdaOut => P(5)(688));
U_G6689: entity G port map(lamdaA => P(6)(673),lamdaB => P(6)(689),s => s(6)(337),lamdaOut => P(5)(689));
U_G6690: entity G port map(lamdaA => P(6)(674),lamdaB => P(6)(690),s => s(6)(338),lamdaOut => P(5)(690));
U_G6691: entity G port map(lamdaA => P(6)(675),lamdaB => P(6)(691),s => s(6)(339),lamdaOut => P(5)(691));
U_G6692: entity G port map(lamdaA => P(6)(676),lamdaB => P(6)(692),s => s(6)(340),lamdaOut => P(5)(692));
U_G6693: entity G port map(lamdaA => P(6)(677),lamdaB => P(6)(693),s => s(6)(341),lamdaOut => P(5)(693));
U_G6694: entity G port map(lamdaA => P(6)(678),lamdaB => P(6)(694),s => s(6)(342),lamdaOut => P(5)(694));
U_G6695: entity G port map(lamdaA => P(6)(679),lamdaB => P(6)(695),s => s(6)(343),lamdaOut => P(5)(695));
U_G6696: entity G port map(lamdaA => P(6)(680),lamdaB => P(6)(696),s => s(6)(344),lamdaOut => P(5)(696));
U_G6697: entity G port map(lamdaA => P(6)(681),lamdaB => P(6)(697),s => s(6)(345),lamdaOut => P(5)(697));
U_G6698: entity G port map(lamdaA => P(6)(682),lamdaB => P(6)(698),s => s(6)(346),lamdaOut => P(5)(698));
U_G6699: entity G port map(lamdaA => P(6)(683),lamdaB => P(6)(699),s => s(6)(347),lamdaOut => P(5)(699));
U_G6700: entity G port map(lamdaA => P(6)(684),lamdaB => P(6)(700),s => s(6)(348),lamdaOut => P(5)(700));
U_G6701: entity G port map(lamdaA => P(6)(685),lamdaB => P(6)(701),s => s(6)(349),lamdaOut => P(5)(701));
U_G6702: entity G port map(lamdaA => P(6)(686),lamdaB => P(6)(702),s => s(6)(350),lamdaOut => P(5)(702));
U_G6703: entity G port map(lamdaA => P(6)(687),lamdaB => P(6)(703),s => s(6)(351),lamdaOut => P(5)(703));
U_F6704: entity F port map(lamdaA => P(6)(704),lamdaB => P(6)(720),lamdaOut => P(5)(704));
U_F6705: entity F port map(lamdaA => P(6)(705),lamdaB => P(6)(721),lamdaOut => P(5)(705));
U_F6706: entity F port map(lamdaA => P(6)(706),lamdaB => P(6)(722),lamdaOut => P(5)(706));
U_F6707: entity F port map(lamdaA => P(6)(707),lamdaB => P(6)(723),lamdaOut => P(5)(707));
U_F6708: entity F port map(lamdaA => P(6)(708),lamdaB => P(6)(724),lamdaOut => P(5)(708));
U_F6709: entity F port map(lamdaA => P(6)(709),lamdaB => P(6)(725),lamdaOut => P(5)(709));
U_F6710: entity F port map(lamdaA => P(6)(710),lamdaB => P(6)(726),lamdaOut => P(5)(710));
U_F6711: entity F port map(lamdaA => P(6)(711),lamdaB => P(6)(727),lamdaOut => P(5)(711));
U_F6712: entity F port map(lamdaA => P(6)(712),lamdaB => P(6)(728),lamdaOut => P(5)(712));
U_F6713: entity F port map(lamdaA => P(6)(713),lamdaB => P(6)(729),lamdaOut => P(5)(713));
U_F6714: entity F port map(lamdaA => P(6)(714),lamdaB => P(6)(730),lamdaOut => P(5)(714));
U_F6715: entity F port map(lamdaA => P(6)(715),lamdaB => P(6)(731),lamdaOut => P(5)(715));
U_F6716: entity F port map(lamdaA => P(6)(716),lamdaB => P(6)(732),lamdaOut => P(5)(716));
U_F6717: entity F port map(lamdaA => P(6)(717),lamdaB => P(6)(733),lamdaOut => P(5)(717));
U_F6718: entity F port map(lamdaA => P(6)(718),lamdaB => P(6)(734),lamdaOut => P(5)(718));
U_F6719: entity F port map(lamdaA => P(6)(719),lamdaB => P(6)(735),lamdaOut => P(5)(719));
U_G6720: entity G port map(lamdaA => P(6)(704),lamdaB => P(6)(720),s => s(6)(352),lamdaOut => P(5)(720));
U_G6721: entity G port map(lamdaA => P(6)(705),lamdaB => P(6)(721),s => s(6)(353),lamdaOut => P(5)(721));
U_G6722: entity G port map(lamdaA => P(6)(706),lamdaB => P(6)(722),s => s(6)(354),lamdaOut => P(5)(722));
U_G6723: entity G port map(lamdaA => P(6)(707),lamdaB => P(6)(723),s => s(6)(355),lamdaOut => P(5)(723));
U_G6724: entity G port map(lamdaA => P(6)(708),lamdaB => P(6)(724),s => s(6)(356),lamdaOut => P(5)(724));
U_G6725: entity G port map(lamdaA => P(6)(709),lamdaB => P(6)(725),s => s(6)(357),lamdaOut => P(5)(725));
U_G6726: entity G port map(lamdaA => P(6)(710),lamdaB => P(6)(726),s => s(6)(358),lamdaOut => P(5)(726));
U_G6727: entity G port map(lamdaA => P(6)(711),lamdaB => P(6)(727),s => s(6)(359),lamdaOut => P(5)(727));
U_G6728: entity G port map(lamdaA => P(6)(712),lamdaB => P(6)(728),s => s(6)(360),lamdaOut => P(5)(728));
U_G6729: entity G port map(lamdaA => P(6)(713),lamdaB => P(6)(729),s => s(6)(361),lamdaOut => P(5)(729));
U_G6730: entity G port map(lamdaA => P(6)(714),lamdaB => P(6)(730),s => s(6)(362),lamdaOut => P(5)(730));
U_G6731: entity G port map(lamdaA => P(6)(715),lamdaB => P(6)(731),s => s(6)(363),lamdaOut => P(5)(731));
U_G6732: entity G port map(lamdaA => P(6)(716),lamdaB => P(6)(732),s => s(6)(364),lamdaOut => P(5)(732));
U_G6733: entity G port map(lamdaA => P(6)(717),lamdaB => P(6)(733),s => s(6)(365),lamdaOut => P(5)(733));
U_G6734: entity G port map(lamdaA => P(6)(718),lamdaB => P(6)(734),s => s(6)(366),lamdaOut => P(5)(734));
U_G6735: entity G port map(lamdaA => P(6)(719),lamdaB => P(6)(735),s => s(6)(367),lamdaOut => P(5)(735));
U_F6736: entity F port map(lamdaA => P(6)(736),lamdaB => P(6)(752),lamdaOut => P(5)(736));
U_F6737: entity F port map(lamdaA => P(6)(737),lamdaB => P(6)(753),lamdaOut => P(5)(737));
U_F6738: entity F port map(lamdaA => P(6)(738),lamdaB => P(6)(754),lamdaOut => P(5)(738));
U_F6739: entity F port map(lamdaA => P(6)(739),lamdaB => P(6)(755),lamdaOut => P(5)(739));
U_F6740: entity F port map(lamdaA => P(6)(740),lamdaB => P(6)(756),lamdaOut => P(5)(740));
U_F6741: entity F port map(lamdaA => P(6)(741),lamdaB => P(6)(757),lamdaOut => P(5)(741));
U_F6742: entity F port map(lamdaA => P(6)(742),lamdaB => P(6)(758),lamdaOut => P(5)(742));
U_F6743: entity F port map(lamdaA => P(6)(743),lamdaB => P(6)(759),lamdaOut => P(5)(743));
U_F6744: entity F port map(lamdaA => P(6)(744),lamdaB => P(6)(760),lamdaOut => P(5)(744));
U_F6745: entity F port map(lamdaA => P(6)(745),lamdaB => P(6)(761),lamdaOut => P(5)(745));
U_F6746: entity F port map(lamdaA => P(6)(746),lamdaB => P(6)(762),lamdaOut => P(5)(746));
U_F6747: entity F port map(lamdaA => P(6)(747),lamdaB => P(6)(763),lamdaOut => P(5)(747));
U_F6748: entity F port map(lamdaA => P(6)(748),lamdaB => P(6)(764),lamdaOut => P(5)(748));
U_F6749: entity F port map(lamdaA => P(6)(749),lamdaB => P(6)(765),lamdaOut => P(5)(749));
U_F6750: entity F port map(lamdaA => P(6)(750),lamdaB => P(6)(766),lamdaOut => P(5)(750));
U_F6751: entity F port map(lamdaA => P(6)(751),lamdaB => P(6)(767),lamdaOut => P(5)(751));
U_G6752: entity G port map(lamdaA => P(6)(736),lamdaB => P(6)(752),s => s(6)(368),lamdaOut => P(5)(752));
U_G6753: entity G port map(lamdaA => P(6)(737),lamdaB => P(6)(753),s => s(6)(369),lamdaOut => P(5)(753));
U_G6754: entity G port map(lamdaA => P(6)(738),lamdaB => P(6)(754),s => s(6)(370),lamdaOut => P(5)(754));
U_G6755: entity G port map(lamdaA => P(6)(739),lamdaB => P(6)(755),s => s(6)(371),lamdaOut => P(5)(755));
U_G6756: entity G port map(lamdaA => P(6)(740),lamdaB => P(6)(756),s => s(6)(372),lamdaOut => P(5)(756));
U_G6757: entity G port map(lamdaA => P(6)(741),lamdaB => P(6)(757),s => s(6)(373),lamdaOut => P(5)(757));
U_G6758: entity G port map(lamdaA => P(6)(742),lamdaB => P(6)(758),s => s(6)(374),lamdaOut => P(5)(758));
U_G6759: entity G port map(lamdaA => P(6)(743),lamdaB => P(6)(759),s => s(6)(375),lamdaOut => P(5)(759));
U_G6760: entity G port map(lamdaA => P(6)(744),lamdaB => P(6)(760),s => s(6)(376),lamdaOut => P(5)(760));
U_G6761: entity G port map(lamdaA => P(6)(745),lamdaB => P(6)(761),s => s(6)(377),lamdaOut => P(5)(761));
U_G6762: entity G port map(lamdaA => P(6)(746),lamdaB => P(6)(762),s => s(6)(378),lamdaOut => P(5)(762));
U_G6763: entity G port map(lamdaA => P(6)(747),lamdaB => P(6)(763),s => s(6)(379),lamdaOut => P(5)(763));
U_G6764: entity G port map(lamdaA => P(6)(748),lamdaB => P(6)(764),s => s(6)(380),lamdaOut => P(5)(764));
U_G6765: entity G port map(lamdaA => P(6)(749),lamdaB => P(6)(765),s => s(6)(381),lamdaOut => P(5)(765));
U_G6766: entity G port map(lamdaA => P(6)(750),lamdaB => P(6)(766),s => s(6)(382),lamdaOut => P(5)(766));
U_G6767: entity G port map(lamdaA => P(6)(751),lamdaB => P(6)(767),s => s(6)(383),lamdaOut => P(5)(767));
U_F6768: entity F port map(lamdaA => P(6)(768),lamdaB => P(6)(784),lamdaOut => P(5)(768));
U_F6769: entity F port map(lamdaA => P(6)(769),lamdaB => P(6)(785),lamdaOut => P(5)(769));
U_F6770: entity F port map(lamdaA => P(6)(770),lamdaB => P(6)(786),lamdaOut => P(5)(770));
U_F6771: entity F port map(lamdaA => P(6)(771),lamdaB => P(6)(787),lamdaOut => P(5)(771));
U_F6772: entity F port map(lamdaA => P(6)(772),lamdaB => P(6)(788),lamdaOut => P(5)(772));
U_F6773: entity F port map(lamdaA => P(6)(773),lamdaB => P(6)(789),lamdaOut => P(5)(773));
U_F6774: entity F port map(lamdaA => P(6)(774),lamdaB => P(6)(790),lamdaOut => P(5)(774));
U_F6775: entity F port map(lamdaA => P(6)(775),lamdaB => P(6)(791),lamdaOut => P(5)(775));
U_F6776: entity F port map(lamdaA => P(6)(776),lamdaB => P(6)(792),lamdaOut => P(5)(776));
U_F6777: entity F port map(lamdaA => P(6)(777),lamdaB => P(6)(793),lamdaOut => P(5)(777));
U_F6778: entity F port map(lamdaA => P(6)(778),lamdaB => P(6)(794),lamdaOut => P(5)(778));
U_F6779: entity F port map(lamdaA => P(6)(779),lamdaB => P(6)(795),lamdaOut => P(5)(779));
U_F6780: entity F port map(lamdaA => P(6)(780),lamdaB => P(6)(796),lamdaOut => P(5)(780));
U_F6781: entity F port map(lamdaA => P(6)(781),lamdaB => P(6)(797),lamdaOut => P(5)(781));
U_F6782: entity F port map(lamdaA => P(6)(782),lamdaB => P(6)(798),lamdaOut => P(5)(782));
U_F6783: entity F port map(lamdaA => P(6)(783),lamdaB => P(6)(799),lamdaOut => P(5)(783));
U_G6784: entity G port map(lamdaA => P(6)(768),lamdaB => P(6)(784),s => s(6)(384),lamdaOut => P(5)(784));
U_G6785: entity G port map(lamdaA => P(6)(769),lamdaB => P(6)(785),s => s(6)(385),lamdaOut => P(5)(785));
U_G6786: entity G port map(lamdaA => P(6)(770),lamdaB => P(6)(786),s => s(6)(386),lamdaOut => P(5)(786));
U_G6787: entity G port map(lamdaA => P(6)(771),lamdaB => P(6)(787),s => s(6)(387),lamdaOut => P(5)(787));
U_G6788: entity G port map(lamdaA => P(6)(772),lamdaB => P(6)(788),s => s(6)(388),lamdaOut => P(5)(788));
U_G6789: entity G port map(lamdaA => P(6)(773),lamdaB => P(6)(789),s => s(6)(389),lamdaOut => P(5)(789));
U_G6790: entity G port map(lamdaA => P(6)(774),lamdaB => P(6)(790),s => s(6)(390),lamdaOut => P(5)(790));
U_G6791: entity G port map(lamdaA => P(6)(775),lamdaB => P(6)(791),s => s(6)(391),lamdaOut => P(5)(791));
U_G6792: entity G port map(lamdaA => P(6)(776),lamdaB => P(6)(792),s => s(6)(392),lamdaOut => P(5)(792));
U_G6793: entity G port map(lamdaA => P(6)(777),lamdaB => P(6)(793),s => s(6)(393),lamdaOut => P(5)(793));
U_G6794: entity G port map(lamdaA => P(6)(778),lamdaB => P(6)(794),s => s(6)(394),lamdaOut => P(5)(794));
U_G6795: entity G port map(lamdaA => P(6)(779),lamdaB => P(6)(795),s => s(6)(395),lamdaOut => P(5)(795));
U_G6796: entity G port map(lamdaA => P(6)(780),lamdaB => P(6)(796),s => s(6)(396),lamdaOut => P(5)(796));
U_G6797: entity G port map(lamdaA => P(6)(781),lamdaB => P(6)(797),s => s(6)(397),lamdaOut => P(5)(797));
U_G6798: entity G port map(lamdaA => P(6)(782),lamdaB => P(6)(798),s => s(6)(398),lamdaOut => P(5)(798));
U_G6799: entity G port map(lamdaA => P(6)(783),lamdaB => P(6)(799),s => s(6)(399),lamdaOut => P(5)(799));
U_F6800: entity F port map(lamdaA => P(6)(800),lamdaB => P(6)(816),lamdaOut => P(5)(800));
U_F6801: entity F port map(lamdaA => P(6)(801),lamdaB => P(6)(817),lamdaOut => P(5)(801));
U_F6802: entity F port map(lamdaA => P(6)(802),lamdaB => P(6)(818),lamdaOut => P(5)(802));
U_F6803: entity F port map(lamdaA => P(6)(803),lamdaB => P(6)(819),lamdaOut => P(5)(803));
U_F6804: entity F port map(lamdaA => P(6)(804),lamdaB => P(6)(820),lamdaOut => P(5)(804));
U_F6805: entity F port map(lamdaA => P(6)(805),lamdaB => P(6)(821),lamdaOut => P(5)(805));
U_F6806: entity F port map(lamdaA => P(6)(806),lamdaB => P(6)(822),lamdaOut => P(5)(806));
U_F6807: entity F port map(lamdaA => P(6)(807),lamdaB => P(6)(823),lamdaOut => P(5)(807));
U_F6808: entity F port map(lamdaA => P(6)(808),lamdaB => P(6)(824),lamdaOut => P(5)(808));
U_F6809: entity F port map(lamdaA => P(6)(809),lamdaB => P(6)(825),lamdaOut => P(5)(809));
U_F6810: entity F port map(lamdaA => P(6)(810),lamdaB => P(6)(826),lamdaOut => P(5)(810));
U_F6811: entity F port map(lamdaA => P(6)(811),lamdaB => P(6)(827),lamdaOut => P(5)(811));
U_F6812: entity F port map(lamdaA => P(6)(812),lamdaB => P(6)(828),lamdaOut => P(5)(812));
U_F6813: entity F port map(lamdaA => P(6)(813),lamdaB => P(6)(829),lamdaOut => P(5)(813));
U_F6814: entity F port map(lamdaA => P(6)(814),lamdaB => P(6)(830),lamdaOut => P(5)(814));
U_F6815: entity F port map(lamdaA => P(6)(815),lamdaB => P(6)(831),lamdaOut => P(5)(815));
U_G6816: entity G port map(lamdaA => P(6)(800),lamdaB => P(6)(816),s => s(6)(400),lamdaOut => P(5)(816));
U_G6817: entity G port map(lamdaA => P(6)(801),lamdaB => P(6)(817),s => s(6)(401),lamdaOut => P(5)(817));
U_G6818: entity G port map(lamdaA => P(6)(802),lamdaB => P(6)(818),s => s(6)(402),lamdaOut => P(5)(818));
U_G6819: entity G port map(lamdaA => P(6)(803),lamdaB => P(6)(819),s => s(6)(403),lamdaOut => P(5)(819));
U_G6820: entity G port map(lamdaA => P(6)(804),lamdaB => P(6)(820),s => s(6)(404),lamdaOut => P(5)(820));
U_G6821: entity G port map(lamdaA => P(6)(805),lamdaB => P(6)(821),s => s(6)(405),lamdaOut => P(5)(821));
U_G6822: entity G port map(lamdaA => P(6)(806),lamdaB => P(6)(822),s => s(6)(406),lamdaOut => P(5)(822));
U_G6823: entity G port map(lamdaA => P(6)(807),lamdaB => P(6)(823),s => s(6)(407),lamdaOut => P(5)(823));
U_G6824: entity G port map(lamdaA => P(6)(808),lamdaB => P(6)(824),s => s(6)(408),lamdaOut => P(5)(824));
U_G6825: entity G port map(lamdaA => P(6)(809),lamdaB => P(6)(825),s => s(6)(409),lamdaOut => P(5)(825));
U_G6826: entity G port map(lamdaA => P(6)(810),lamdaB => P(6)(826),s => s(6)(410),lamdaOut => P(5)(826));
U_G6827: entity G port map(lamdaA => P(6)(811),lamdaB => P(6)(827),s => s(6)(411),lamdaOut => P(5)(827));
U_G6828: entity G port map(lamdaA => P(6)(812),lamdaB => P(6)(828),s => s(6)(412),lamdaOut => P(5)(828));
U_G6829: entity G port map(lamdaA => P(6)(813),lamdaB => P(6)(829),s => s(6)(413),lamdaOut => P(5)(829));
U_G6830: entity G port map(lamdaA => P(6)(814),lamdaB => P(6)(830),s => s(6)(414),lamdaOut => P(5)(830));
U_G6831: entity G port map(lamdaA => P(6)(815),lamdaB => P(6)(831),s => s(6)(415),lamdaOut => P(5)(831));
U_F6832: entity F port map(lamdaA => P(6)(832),lamdaB => P(6)(848),lamdaOut => P(5)(832));
U_F6833: entity F port map(lamdaA => P(6)(833),lamdaB => P(6)(849),lamdaOut => P(5)(833));
U_F6834: entity F port map(lamdaA => P(6)(834),lamdaB => P(6)(850),lamdaOut => P(5)(834));
U_F6835: entity F port map(lamdaA => P(6)(835),lamdaB => P(6)(851),lamdaOut => P(5)(835));
U_F6836: entity F port map(lamdaA => P(6)(836),lamdaB => P(6)(852),lamdaOut => P(5)(836));
U_F6837: entity F port map(lamdaA => P(6)(837),lamdaB => P(6)(853),lamdaOut => P(5)(837));
U_F6838: entity F port map(lamdaA => P(6)(838),lamdaB => P(6)(854),lamdaOut => P(5)(838));
U_F6839: entity F port map(lamdaA => P(6)(839),lamdaB => P(6)(855),lamdaOut => P(5)(839));
U_F6840: entity F port map(lamdaA => P(6)(840),lamdaB => P(6)(856),lamdaOut => P(5)(840));
U_F6841: entity F port map(lamdaA => P(6)(841),lamdaB => P(6)(857),lamdaOut => P(5)(841));
U_F6842: entity F port map(lamdaA => P(6)(842),lamdaB => P(6)(858),lamdaOut => P(5)(842));
U_F6843: entity F port map(lamdaA => P(6)(843),lamdaB => P(6)(859),lamdaOut => P(5)(843));
U_F6844: entity F port map(lamdaA => P(6)(844),lamdaB => P(6)(860),lamdaOut => P(5)(844));
U_F6845: entity F port map(lamdaA => P(6)(845),lamdaB => P(6)(861),lamdaOut => P(5)(845));
U_F6846: entity F port map(lamdaA => P(6)(846),lamdaB => P(6)(862),lamdaOut => P(5)(846));
U_F6847: entity F port map(lamdaA => P(6)(847),lamdaB => P(6)(863),lamdaOut => P(5)(847));
U_G6848: entity G port map(lamdaA => P(6)(832),lamdaB => P(6)(848),s => s(6)(416),lamdaOut => P(5)(848));
U_G6849: entity G port map(lamdaA => P(6)(833),lamdaB => P(6)(849),s => s(6)(417),lamdaOut => P(5)(849));
U_G6850: entity G port map(lamdaA => P(6)(834),lamdaB => P(6)(850),s => s(6)(418),lamdaOut => P(5)(850));
U_G6851: entity G port map(lamdaA => P(6)(835),lamdaB => P(6)(851),s => s(6)(419),lamdaOut => P(5)(851));
U_G6852: entity G port map(lamdaA => P(6)(836),lamdaB => P(6)(852),s => s(6)(420),lamdaOut => P(5)(852));
U_G6853: entity G port map(lamdaA => P(6)(837),lamdaB => P(6)(853),s => s(6)(421),lamdaOut => P(5)(853));
U_G6854: entity G port map(lamdaA => P(6)(838),lamdaB => P(6)(854),s => s(6)(422),lamdaOut => P(5)(854));
U_G6855: entity G port map(lamdaA => P(6)(839),lamdaB => P(6)(855),s => s(6)(423),lamdaOut => P(5)(855));
U_G6856: entity G port map(lamdaA => P(6)(840),lamdaB => P(6)(856),s => s(6)(424),lamdaOut => P(5)(856));
U_G6857: entity G port map(lamdaA => P(6)(841),lamdaB => P(6)(857),s => s(6)(425),lamdaOut => P(5)(857));
U_G6858: entity G port map(lamdaA => P(6)(842),lamdaB => P(6)(858),s => s(6)(426),lamdaOut => P(5)(858));
U_G6859: entity G port map(lamdaA => P(6)(843),lamdaB => P(6)(859),s => s(6)(427),lamdaOut => P(5)(859));
U_G6860: entity G port map(lamdaA => P(6)(844),lamdaB => P(6)(860),s => s(6)(428),lamdaOut => P(5)(860));
U_G6861: entity G port map(lamdaA => P(6)(845),lamdaB => P(6)(861),s => s(6)(429),lamdaOut => P(5)(861));
U_G6862: entity G port map(lamdaA => P(6)(846),lamdaB => P(6)(862),s => s(6)(430),lamdaOut => P(5)(862));
U_G6863: entity G port map(lamdaA => P(6)(847),lamdaB => P(6)(863),s => s(6)(431),lamdaOut => P(5)(863));
U_F6864: entity F port map(lamdaA => P(6)(864),lamdaB => P(6)(880),lamdaOut => P(5)(864));
U_F6865: entity F port map(lamdaA => P(6)(865),lamdaB => P(6)(881),lamdaOut => P(5)(865));
U_F6866: entity F port map(lamdaA => P(6)(866),lamdaB => P(6)(882),lamdaOut => P(5)(866));
U_F6867: entity F port map(lamdaA => P(6)(867),lamdaB => P(6)(883),lamdaOut => P(5)(867));
U_F6868: entity F port map(lamdaA => P(6)(868),lamdaB => P(6)(884),lamdaOut => P(5)(868));
U_F6869: entity F port map(lamdaA => P(6)(869),lamdaB => P(6)(885),lamdaOut => P(5)(869));
U_F6870: entity F port map(lamdaA => P(6)(870),lamdaB => P(6)(886),lamdaOut => P(5)(870));
U_F6871: entity F port map(lamdaA => P(6)(871),lamdaB => P(6)(887),lamdaOut => P(5)(871));
U_F6872: entity F port map(lamdaA => P(6)(872),lamdaB => P(6)(888),lamdaOut => P(5)(872));
U_F6873: entity F port map(lamdaA => P(6)(873),lamdaB => P(6)(889),lamdaOut => P(5)(873));
U_F6874: entity F port map(lamdaA => P(6)(874),lamdaB => P(6)(890),lamdaOut => P(5)(874));
U_F6875: entity F port map(lamdaA => P(6)(875),lamdaB => P(6)(891),lamdaOut => P(5)(875));
U_F6876: entity F port map(lamdaA => P(6)(876),lamdaB => P(6)(892),lamdaOut => P(5)(876));
U_F6877: entity F port map(lamdaA => P(6)(877),lamdaB => P(6)(893),lamdaOut => P(5)(877));
U_F6878: entity F port map(lamdaA => P(6)(878),lamdaB => P(6)(894),lamdaOut => P(5)(878));
U_F6879: entity F port map(lamdaA => P(6)(879),lamdaB => P(6)(895),lamdaOut => P(5)(879));
U_G6880: entity G port map(lamdaA => P(6)(864),lamdaB => P(6)(880),s => s(6)(432),lamdaOut => P(5)(880));
U_G6881: entity G port map(lamdaA => P(6)(865),lamdaB => P(6)(881),s => s(6)(433),lamdaOut => P(5)(881));
U_G6882: entity G port map(lamdaA => P(6)(866),lamdaB => P(6)(882),s => s(6)(434),lamdaOut => P(5)(882));
U_G6883: entity G port map(lamdaA => P(6)(867),lamdaB => P(6)(883),s => s(6)(435),lamdaOut => P(5)(883));
U_G6884: entity G port map(lamdaA => P(6)(868),lamdaB => P(6)(884),s => s(6)(436),lamdaOut => P(5)(884));
U_G6885: entity G port map(lamdaA => P(6)(869),lamdaB => P(6)(885),s => s(6)(437),lamdaOut => P(5)(885));
U_G6886: entity G port map(lamdaA => P(6)(870),lamdaB => P(6)(886),s => s(6)(438),lamdaOut => P(5)(886));
U_G6887: entity G port map(lamdaA => P(6)(871),lamdaB => P(6)(887),s => s(6)(439),lamdaOut => P(5)(887));
U_G6888: entity G port map(lamdaA => P(6)(872),lamdaB => P(6)(888),s => s(6)(440),lamdaOut => P(5)(888));
U_G6889: entity G port map(lamdaA => P(6)(873),lamdaB => P(6)(889),s => s(6)(441),lamdaOut => P(5)(889));
U_G6890: entity G port map(lamdaA => P(6)(874),lamdaB => P(6)(890),s => s(6)(442),lamdaOut => P(5)(890));
U_G6891: entity G port map(lamdaA => P(6)(875),lamdaB => P(6)(891),s => s(6)(443),lamdaOut => P(5)(891));
U_G6892: entity G port map(lamdaA => P(6)(876),lamdaB => P(6)(892),s => s(6)(444),lamdaOut => P(5)(892));
U_G6893: entity G port map(lamdaA => P(6)(877),lamdaB => P(6)(893),s => s(6)(445),lamdaOut => P(5)(893));
U_G6894: entity G port map(lamdaA => P(6)(878),lamdaB => P(6)(894),s => s(6)(446),lamdaOut => P(5)(894));
U_G6895: entity G port map(lamdaA => P(6)(879),lamdaB => P(6)(895),s => s(6)(447),lamdaOut => P(5)(895));
U_F6896: entity F port map(lamdaA => P(6)(896),lamdaB => P(6)(912),lamdaOut => P(5)(896));
U_F6897: entity F port map(lamdaA => P(6)(897),lamdaB => P(6)(913),lamdaOut => P(5)(897));
U_F6898: entity F port map(lamdaA => P(6)(898),lamdaB => P(6)(914),lamdaOut => P(5)(898));
U_F6899: entity F port map(lamdaA => P(6)(899),lamdaB => P(6)(915),lamdaOut => P(5)(899));
U_F6900: entity F port map(lamdaA => P(6)(900),lamdaB => P(6)(916),lamdaOut => P(5)(900));
U_F6901: entity F port map(lamdaA => P(6)(901),lamdaB => P(6)(917),lamdaOut => P(5)(901));
U_F6902: entity F port map(lamdaA => P(6)(902),lamdaB => P(6)(918),lamdaOut => P(5)(902));
U_F6903: entity F port map(lamdaA => P(6)(903),lamdaB => P(6)(919),lamdaOut => P(5)(903));
U_F6904: entity F port map(lamdaA => P(6)(904),lamdaB => P(6)(920),lamdaOut => P(5)(904));
U_F6905: entity F port map(lamdaA => P(6)(905),lamdaB => P(6)(921),lamdaOut => P(5)(905));
U_F6906: entity F port map(lamdaA => P(6)(906),lamdaB => P(6)(922),lamdaOut => P(5)(906));
U_F6907: entity F port map(lamdaA => P(6)(907),lamdaB => P(6)(923),lamdaOut => P(5)(907));
U_F6908: entity F port map(lamdaA => P(6)(908),lamdaB => P(6)(924),lamdaOut => P(5)(908));
U_F6909: entity F port map(lamdaA => P(6)(909),lamdaB => P(6)(925),lamdaOut => P(5)(909));
U_F6910: entity F port map(lamdaA => P(6)(910),lamdaB => P(6)(926),lamdaOut => P(5)(910));
U_F6911: entity F port map(lamdaA => P(6)(911),lamdaB => P(6)(927),lamdaOut => P(5)(911));
U_G6912: entity G port map(lamdaA => P(6)(896),lamdaB => P(6)(912),s => s(6)(448),lamdaOut => P(5)(912));
U_G6913: entity G port map(lamdaA => P(6)(897),lamdaB => P(6)(913),s => s(6)(449),lamdaOut => P(5)(913));
U_G6914: entity G port map(lamdaA => P(6)(898),lamdaB => P(6)(914),s => s(6)(450),lamdaOut => P(5)(914));
U_G6915: entity G port map(lamdaA => P(6)(899),lamdaB => P(6)(915),s => s(6)(451),lamdaOut => P(5)(915));
U_G6916: entity G port map(lamdaA => P(6)(900),lamdaB => P(6)(916),s => s(6)(452),lamdaOut => P(5)(916));
U_G6917: entity G port map(lamdaA => P(6)(901),lamdaB => P(6)(917),s => s(6)(453),lamdaOut => P(5)(917));
U_G6918: entity G port map(lamdaA => P(6)(902),lamdaB => P(6)(918),s => s(6)(454),lamdaOut => P(5)(918));
U_G6919: entity G port map(lamdaA => P(6)(903),lamdaB => P(6)(919),s => s(6)(455),lamdaOut => P(5)(919));
U_G6920: entity G port map(lamdaA => P(6)(904),lamdaB => P(6)(920),s => s(6)(456),lamdaOut => P(5)(920));
U_G6921: entity G port map(lamdaA => P(6)(905),lamdaB => P(6)(921),s => s(6)(457),lamdaOut => P(5)(921));
U_G6922: entity G port map(lamdaA => P(6)(906),lamdaB => P(6)(922),s => s(6)(458),lamdaOut => P(5)(922));
U_G6923: entity G port map(lamdaA => P(6)(907),lamdaB => P(6)(923),s => s(6)(459),lamdaOut => P(5)(923));
U_G6924: entity G port map(lamdaA => P(6)(908),lamdaB => P(6)(924),s => s(6)(460),lamdaOut => P(5)(924));
U_G6925: entity G port map(lamdaA => P(6)(909),lamdaB => P(6)(925),s => s(6)(461),lamdaOut => P(5)(925));
U_G6926: entity G port map(lamdaA => P(6)(910),lamdaB => P(6)(926),s => s(6)(462),lamdaOut => P(5)(926));
U_G6927: entity G port map(lamdaA => P(6)(911),lamdaB => P(6)(927),s => s(6)(463),lamdaOut => P(5)(927));
U_F6928: entity F port map(lamdaA => P(6)(928),lamdaB => P(6)(944),lamdaOut => P(5)(928));
U_F6929: entity F port map(lamdaA => P(6)(929),lamdaB => P(6)(945),lamdaOut => P(5)(929));
U_F6930: entity F port map(lamdaA => P(6)(930),lamdaB => P(6)(946),lamdaOut => P(5)(930));
U_F6931: entity F port map(lamdaA => P(6)(931),lamdaB => P(6)(947),lamdaOut => P(5)(931));
U_F6932: entity F port map(lamdaA => P(6)(932),lamdaB => P(6)(948),lamdaOut => P(5)(932));
U_F6933: entity F port map(lamdaA => P(6)(933),lamdaB => P(6)(949),lamdaOut => P(5)(933));
U_F6934: entity F port map(lamdaA => P(6)(934),lamdaB => P(6)(950),lamdaOut => P(5)(934));
U_F6935: entity F port map(lamdaA => P(6)(935),lamdaB => P(6)(951),lamdaOut => P(5)(935));
U_F6936: entity F port map(lamdaA => P(6)(936),lamdaB => P(6)(952),lamdaOut => P(5)(936));
U_F6937: entity F port map(lamdaA => P(6)(937),lamdaB => P(6)(953),lamdaOut => P(5)(937));
U_F6938: entity F port map(lamdaA => P(6)(938),lamdaB => P(6)(954),lamdaOut => P(5)(938));
U_F6939: entity F port map(lamdaA => P(6)(939),lamdaB => P(6)(955),lamdaOut => P(5)(939));
U_F6940: entity F port map(lamdaA => P(6)(940),lamdaB => P(6)(956),lamdaOut => P(5)(940));
U_F6941: entity F port map(lamdaA => P(6)(941),lamdaB => P(6)(957),lamdaOut => P(5)(941));
U_F6942: entity F port map(lamdaA => P(6)(942),lamdaB => P(6)(958),lamdaOut => P(5)(942));
U_F6943: entity F port map(lamdaA => P(6)(943),lamdaB => P(6)(959),lamdaOut => P(5)(943));
U_G6944: entity G port map(lamdaA => P(6)(928),lamdaB => P(6)(944),s => s(6)(464),lamdaOut => P(5)(944));
U_G6945: entity G port map(lamdaA => P(6)(929),lamdaB => P(6)(945),s => s(6)(465),lamdaOut => P(5)(945));
U_G6946: entity G port map(lamdaA => P(6)(930),lamdaB => P(6)(946),s => s(6)(466),lamdaOut => P(5)(946));
U_G6947: entity G port map(lamdaA => P(6)(931),lamdaB => P(6)(947),s => s(6)(467),lamdaOut => P(5)(947));
U_G6948: entity G port map(lamdaA => P(6)(932),lamdaB => P(6)(948),s => s(6)(468),lamdaOut => P(5)(948));
U_G6949: entity G port map(lamdaA => P(6)(933),lamdaB => P(6)(949),s => s(6)(469),lamdaOut => P(5)(949));
U_G6950: entity G port map(lamdaA => P(6)(934),lamdaB => P(6)(950),s => s(6)(470),lamdaOut => P(5)(950));
U_G6951: entity G port map(lamdaA => P(6)(935),lamdaB => P(6)(951),s => s(6)(471),lamdaOut => P(5)(951));
U_G6952: entity G port map(lamdaA => P(6)(936),lamdaB => P(6)(952),s => s(6)(472),lamdaOut => P(5)(952));
U_G6953: entity G port map(lamdaA => P(6)(937),lamdaB => P(6)(953),s => s(6)(473),lamdaOut => P(5)(953));
U_G6954: entity G port map(lamdaA => P(6)(938),lamdaB => P(6)(954),s => s(6)(474),lamdaOut => P(5)(954));
U_G6955: entity G port map(lamdaA => P(6)(939),lamdaB => P(6)(955),s => s(6)(475),lamdaOut => P(5)(955));
U_G6956: entity G port map(lamdaA => P(6)(940),lamdaB => P(6)(956),s => s(6)(476),lamdaOut => P(5)(956));
U_G6957: entity G port map(lamdaA => P(6)(941),lamdaB => P(6)(957),s => s(6)(477),lamdaOut => P(5)(957));
U_G6958: entity G port map(lamdaA => P(6)(942),lamdaB => P(6)(958),s => s(6)(478),lamdaOut => P(5)(958));
U_G6959: entity G port map(lamdaA => P(6)(943),lamdaB => P(6)(959),s => s(6)(479),lamdaOut => P(5)(959));
U_F6960: entity F port map(lamdaA => P(6)(960),lamdaB => P(6)(976),lamdaOut => P(5)(960));
U_F6961: entity F port map(lamdaA => P(6)(961),lamdaB => P(6)(977),lamdaOut => P(5)(961));
U_F6962: entity F port map(lamdaA => P(6)(962),lamdaB => P(6)(978),lamdaOut => P(5)(962));
U_F6963: entity F port map(lamdaA => P(6)(963),lamdaB => P(6)(979),lamdaOut => P(5)(963));
U_F6964: entity F port map(lamdaA => P(6)(964),lamdaB => P(6)(980),lamdaOut => P(5)(964));
U_F6965: entity F port map(lamdaA => P(6)(965),lamdaB => P(6)(981),lamdaOut => P(5)(965));
U_F6966: entity F port map(lamdaA => P(6)(966),lamdaB => P(6)(982),lamdaOut => P(5)(966));
U_F6967: entity F port map(lamdaA => P(6)(967),lamdaB => P(6)(983),lamdaOut => P(5)(967));
U_F6968: entity F port map(lamdaA => P(6)(968),lamdaB => P(6)(984),lamdaOut => P(5)(968));
U_F6969: entity F port map(lamdaA => P(6)(969),lamdaB => P(6)(985),lamdaOut => P(5)(969));
U_F6970: entity F port map(lamdaA => P(6)(970),lamdaB => P(6)(986),lamdaOut => P(5)(970));
U_F6971: entity F port map(lamdaA => P(6)(971),lamdaB => P(6)(987),lamdaOut => P(5)(971));
U_F6972: entity F port map(lamdaA => P(6)(972),lamdaB => P(6)(988),lamdaOut => P(5)(972));
U_F6973: entity F port map(lamdaA => P(6)(973),lamdaB => P(6)(989),lamdaOut => P(5)(973));
U_F6974: entity F port map(lamdaA => P(6)(974),lamdaB => P(6)(990),lamdaOut => P(5)(974));
U_F6975: entity F port map(lamdaA => P(6)(975),lamdaB => P(6)(991),lamdaOut => P(5)(975));
U_G6976: entity G port map(lamdaA => P(6)(960),lamdaB => P(6)(976),s => s(6)(480),lamdaOut => P(5)(976));
U_G6977: entity G port map(lamdaA => P(6)(961),lamdaB => P(6)(977),s => s(6)(481),lamdaOut => P(5)(977));
U_G6978: entity G port map(lamdaA => P(6)(962),lamdaB => P(6)(978),s => s(6)(482),lamdaOut => P(5)(978));
U_G6979: entity G port map(lamdaA => P(6)(963),lamdaB => P(6)(979),s => s(6)(483),lamdaOut => P(5)(979));
U_G6980: entity G port map(lamdaA => P(6)(964),lamdaB => P(6)(980),s => s(6)(484),lamdaOut => P(5)(980));
U_G6981: entity G port map(lamdaA => P(6)(965),lamdaB => P(6)(981),s => s(6)(485),lamdaOut => P(5)(981));
U_G6982: entity G port map(lamdaA => P(6)(966),lamdaB => P(6)(982),s => s(6)(486),lamdaOut => P(5)(982));
U_G6983: entity G port map(lamdaA => P(6)(967),lamdaB => P(6)(983),s => s(6)(487),lamdaOut => P(5)(983));
U_G6984: entity G port map(lamdaA => P(6)(968),lamdaB => P(6)(984),s => s(6)(488),lamdaOut => P(5)(984));
U_G6985: entity G port map(lamdaA => P(6)(969),lamdaB => P(6)(985),s => s(6)(489),lamdaOut => P(5)(985));
U_G6986: entity G port map(lamdaA => P(6)(970),lamdaB => P(6)(986),s => s(6)(490),lamdaOut => P(5)(986));
U_G6987: entity G port map(lamdaA => P(6)(971),lamdaB => P(6)(987),s => s(6)(491),lamdaOut => P(5)(987));
U_G6988: entity G port map(lamdaA => P(6)(972),lamdaB => P(6)(988),s => s(6)(492),lamdaOut => P(5)(988));
U_G6989: entity G port map(lamdaA => P(6)(973),lamdaB => P(6)(989),s => s(6)(493),lamdaOut => P(5)(989));
U_G6990: entity G port map(lamdaA => P(6)(974),lamdaB => P(6)(990),s => s(6)(494),lamdaOut => P(5)(990));
U_G6991: entity G port map(lamdaA => P(6)(975),lamdaB => P(6)(991),s => s(6)(495),lamdaOut => P(5)(991));
U_F6992: entity F port map(lamdaA => P(6)(992),lamdaB => P(6)(1008),lamdaOut => P(5)(992));
U_F6993: entity F port map(lamdaA => P(6)(993),lamdaB => P(6)(1009),lamdaOut => P(5)(993));
U_F6994: entity F port map(lamdaA => P(6)(994),lamdaB => P(6)(1010),lamdaOut => P(5)(994));
U_F6995: entity F port map(lamdaA => P(6)(995),lamdaB => P(6)(1011),lamdaOut => P(5)(995));
U_F6996: entity F port map(lamdaA => P(6)(996),lamdaB => P(6)(1012),lamdaOut => P(5)(996));
U_F6997: entity F port map(lamdaA => P(6)(997),lamdaB => P(6)(1013),lamdaOut => P(5)(997));
U_F6998: entity F port map(lamdaA => P(6)(998),lamdaB => P(6)(1014),lamdaOut => P(5)(998));
U_F6999: entity F port map(lamdaA => P(6)(999),lamdaB => P(6)(1015),lamdaOut => P(5)(999));
U_F61000: entity F port map(lamdaA => P(6)(1000),lamdaB => P(6)(1016),lamdaOut => P(5)(1000));
U_F61001: entity F port map(lamdaA => P(6)(1001),lamdaB => P(6)(1017),lamdaOut => P(5)(1001));
U_F61002: entity F port map(lamdaA => P(6)(1002),lamdaB => P(6)(1018),lamdaOut => P(5)(1002));
U_F61003: entity F port map(lamdaA => P(6)(1003),lamdaB => P(6)(1019),lamdaOut => P(5)(1003));
U_F61004: entity F port map(lamdaA => P(6)(1004),lamdaB => P(6)(1020),lamdaOut => P(5)(1004));
U_F61005: entity F port map(lamdaA => P(6)(1005),lamdaB => P(6)(1021),lamdaOut => P(5)(1005));
U_F61006: entity F port map(lamdaA => P(6)(1006),lamdaB => P(6)(1022),lamdaOut => P(5)(1006));
U_F61007: entity F port map(lamdaA => P(6)(1007),lamdaB => P(6)(1023),lamdaOut => P(5)(1007));
U_G61008: entity G port map(lamdaA => P(6)(992),lamdaB => P(6)(1008),s => s(6)(496),lamdaOut => P(5)(1008));
U_G61009: entity G port map(lamdaA => P(6)(993),lamdaB => P(6)(1009),s => s(6)(497),lamdaOut => P(5)(1009));
U_G61010: entity G port map(lamdaA => P(6)(994),lamdaB => P(6)(1010),s => s(6)(498),lamdaOut => P(5)(1010));
U_G61011: entity G port map(lamdaA => P(6)(995),lamdaB => P(6)(1011),s => s(6)(499),lamdaOut => P(5)(1011));
U_G61012: entity G port map(lamdaA => P(6)(996),lamdaB => P(6)(1012),s => s(6)(500),lamdaOut => P(5)(1012));
U_G61013: entity G port map(lamdaA => P(6)(997),lamdaB => P(6)(1013),s => s(6)(501),lamdaOut => P(5)(1013));
U_G61014: entity G port map(lamdaA => P(6)(998),lamdaB => P(6)(1014),s => s(6)(502),lamdaOut => P(5)(1014));
U_G61015: entity G port map(lamdaA => P(6)(999),lamdaB => P(6)(1015),s => s(6)(503),lamdaOut => P(5)(1015));
U_G61016: entity G port map(lamdaA => P(6)(1000),lamdaB => P(6)(1016),s => s(6)(504),lamdaOut => P(5)(1016));
U_G61017: entity G port map(lamdaA => P(6)(1001),lamdaB => P(6)(1017),s => s(6)(505),lamdaOut => P(5)(1017));
U_G61018: entity G port map(lamdaA => P(6)(1002),lamdaB => P(6)(1018),s => s(6)(506),lamdaOut => P(5)(1018));
U_G61019: entity G port map(lamdaA => P(6)(1003),lamdaB => P(6)(1019),s => s(6)(507),lamdaOut => P(5)(1019));
U_G61020: entity G port map(lamdaA => P(6)(1004),lamdaB => P(6)(1020),s => s(6)(508),lamdaOut => P(5)(1020));
U_G61021: entity G port map(lamdaA => P(6)(1005),lamdaB => P(6)(1021),s => s(6)(509),lamdaOut => P(5)(1021));
U_G61022: entity G port map(lamdaA => P(6)(1006),lamdaB => P(6)(1022),s => s(6)(510),lamdaOut => P(5)(1022));
U_G61023: entity G port map(lamdaA => P(6)(1007),lamdaB => P(6)(1023),s => s(6)(511),lamdaOut => P(5)(1023));
-- STAGE 4
U_F50: entity F port map(lamdaA => P(5)(0),lamdaB => P(5)(32),lamdaOut => P(4)(0));
U_F51: entity F port map(lamdaA => P(5)(1),lamdaB => P(5)(33),lamdaOut => P(4)(1));
U_F52: entity F port map(lamdaA => P(5)(2),lamdaB => P(5)(34),lamdaOut => P(4)(2));
U_F53: entity F port map(lamdaA => P(5)(3),lamdaB => P(5)(35),lamdaOut => P(4)(3));
U_F54: entity F port map(lamdaA => P(5)(4),lamdaB => P(5)(36),lamdaOut => P(4)(4));
U_F55: entity F port map(lamdaA => P(5)(5),lamdaB => P(5)(37),lamdaOut => P(4)(5));
U_F56: entity F port map(lamdaA => P(5)(6),lamdaB => P(5)(38),lamdaOut => P(4)(6));
U_F57: entity F port map(lamdaA => P(5)(7),lamdaB => P(5)(39),lamdaOut => P(4)(7));
U_F58: entity F port map(lamdaA => P(5)(8),lamdaB => P(5)(40),lamdaOut => P(4)(8));
U_F59: entity F port map(lamdaA => P(5)(9),lamdaB => P(5)(41),lamdaOut => P(4)(9));
U_F510: entity F port map(lamdaA => P(5)(10),lamdaB => P(5)(42),lamdaOut => P(4)(10));
U_F511: entity F port map(lamdaA => P(5)(11),lamdaB => P(5)(43),lamdaOut => P(4)(11));
U_F512: entity F port map(lamdaA => P(5)(12),lamdaB => P(5)(44),lamdaOut => P(4)(12));
U_F513: entity F port map(lamdaA => P(5)(13),lamdaB => P(5)(45),lamdaOut => P(4)(13));
U_F514: entity F port map(lamdaA => P(5)(14),lamdaB => P(5)(46),lamdaOut => P(4)(14));
U_F515: entity F port map(lamdaA => P(5)(15),lamdaB => P(5)(47),lamdaOut => P(4)(15));
U_F516: entity F port map(lamdaA => P(5)(16),lamdaB => P(5)(48),lamdaOut => P(4)(16));
U_F517: entity F port map(lamdaA => P(5)(17),lamdaB => P(5)(49),lamdaOut => P(4)(17));
U_F518: entity F port map(lamdaA => P(5)(18),lamdaB => P(5)(50),lamdaOut => P(4)(18));
U_F519: entity F port map(lamdaA => P(5)(19),lamdaB => P(5)(51),lamdaOut => P(4)(19));
U_F520: entity F port map(lamdaA => P(5)(20),lamdaB => P(5)(52),lamdaOut => P(4)(20));
U_F521: entity F port map(lamdaA => P(5)(21),lamdaB => P(5)(53),lamdaOut => P(4)(21));
U_F522: entity F port map(lamdaA => P(5)(22),lamdaB => P(5)(54),lamdaOut => P(4)(22));
U_F523: entity F port map(lamdaA => P(5)(23),lamdaB => P(5)(55),lamdaOut => P(4)(23));
U_F524: entity F port map(lamdaA => P(5)(24),lamdaB => P(5)(56),lamdaOut => P(4)(24));
U_F525: entity F port map(lamdaA => P(5)(25),lamdaB => P(5)(57),lamdaOut => P(4)(25));
U_F526: entity F port map(lamdaA => P(5)(26),lamdaB => P(5)(58),lamdaOut => P(4)(26));
U_F527: entity F port map(lamdaA => P(5)(27),lamdaB => P(5)(59),lamdaOut => P(4)(27));
U_F528: entity F port map(lamdaA => P(5)(28),lamdaB => P(5)(60),lamdaOut => P(4)(28));
U_F529: entity F port map(lamdaA => P(5)(29),lamdaB => P(5)(61),lamdaOut => P(4)(29));
U_F530: entity F port map(lamdaA => P(5)(30),lamdaB => P(5)(62),lamdaOut => P(4)(30));
U_F531: entity F port map(lamdaA => P(5)(31),lamdaB => P(5)(63),lamdaOut => P(4)(31));
U_G532: entity G port map(lamdaA => P(5)(0),lamdaB => P(5)(32),s => s(5)(0),lamdaOut => P(4)(32));
U_G533: entity G port map(lamdaA => P(5)(1),lamdaB => P(5)(33),s => s(5)(1),lamdaOut => P(4)(33));
U_G534: entity G port map(lamdaA => P(5)(2),lamdaB => P(5)(34),s => s(5)(2),lamdaOut => P(4)(34));
U_G535: entity G port map(lamdaA => P(5)(3),lamdaB => P(5)(35),s => s(5)(3),lamdaOut => P(4)(35));
U_G536: entity G port map(lamdaA => P(5)(4),lamdaB => P(5)(36),s => s(5)(4),lamdaOut => P(4)(36));
U_G537: entity G port map(lamdaA => P(5)(5),lamdaB => P(5)(37),s => s(5)(5),lamdaOut => P(4)(37));
U_G538: entity G port map(lamdaA => P(5)(6),lamdaB => P(5)(38),s => s(5)(6),lamdaOut => P(4)(38));
U_G539: entity G port map(lamdaA => P(5)(7),lamdaB => P(5)(39),s => s(5)(7),lamdaOut => P(4)(39));
U_G540: entity G port map(lamdaA => P(5)(8),lamdaB => P(5)(40),s => s(5)(8),lamdaOut => P(4)(40));
U_G541: entity G port map(lamdaA => P(5)(9),lamdaB => P(5)(41),s => s(5)(9),lamdaOut => P(4)(41));
U_G542: entity G port map(lamdaA => P(5)(10),lamdaB => P(5)(42),s => s(5)(10),lamdaOut => P(4)(42));
U_G543: entity G port map(lamdaA => P(5)(11),lamdaB => P(5)(43),s => s(5)(11),lamdaOut => P(4)(43));
U_G544: entity G port map(lamdaA => P(5)(12),lamdaB => P(5)(44),s => s(5)(12),lamdaOut => P(4)(44));
U_G545: entity G port map(lamdaA => P(5)(13),lamdaB => P(5)(45),s => s(5)(13),lamdaOut => P(4)(45));
U_G546: entity G port map(lamdaA => P(5)(14),lamdaB => P(5)(46),s => s(5)(14),lamdaOut => P(4)(46));
U_G547: entity G port map(lamdaA => P(5)(15),lamdaB => P(5)(47),s => s(5)(15),lamdaOut => P(4)(47));
U_G548: entity G port map(lamdaA => P(5)(16),lamdaB => P(5)(48),s => s(5)(16),lamdaOut => P(4)(48));
U_G549: entity G port map(lamdaA => P(5)(17),lamdaB => P(5)(49),s => s(5)(17),lamdaOut => P(4)(49));
U_G550: entity G port map(lamdaA => P(5)(18),lamdaB => P(5)(50),s => s(5)(18),lamdaOut => P(4)(50));
U_G551: entity G port map(lamdaA => P(5)(19),lamdaB => P(5)(51),s => s(5)(19),lamdaOut => P(4)(51));
U_G552: entity G port map(lamdaA => P(5)(20),lamdaB => P(5)(52),s => s(5)(20),lamdaOut => P(4)(52));
U_G553: entity G port map(lamdaA => P(5)(21),lamdaB => P(5)(53),s => s(5)(21),lamdaOut => P(4)(53));
U_G554: entity G port map(lamdaA => P(5)(22),lamdaB => P(5)(54),s => s(5)(22),lamdaOut => P(4)(54));
U_G555: entity G port map(lamdaA => P(5)(23),lamdaB => P(5)(55),s => s(5)(23),lamdaOut => P(4)(55));
U_G556: entity G port map(lamdaA => P(5)(24),lamdaB => P(5)(56),s => s(5)(24),lamdaOut => P(4)(56));
U_G557: entity G port map(lamdaA => P(5)(25),lamdaB => P(5)(57),s => s(5)(25),lamdaOut => P(4)(57));
U_G558: entity G port map(lamdaA => P(5)(26),lamdaB => P(5)(58),s => s(5)(26),lamdaOut => P(4)(58));
U_G559: entity G port map(lamdaA => P(5)(27),lamdaB => P(5)(59),s => s(5)(27),lamdaOut => P(4)(59));
U_G560: entity G port map(lamdaA => P(5)(28),lamdaB => P(5)(60),s => s(5)(28),lamdaOut => P(4)(60));
U_G561: entity G port map(lamdaA => P(5)(29),lamdaB => P(5)(61),s => s(5)(29),lamdaOut => P(4)(61));
U_G562: entity G port map(lamdaA => P(5)(30),lamdaB => P(5)(62),s => s(5)(30),lamdaOut => P(4)(62));
U_G563: entity G port map(lamdaA => P(5)(31),lamdaB => P(5)(63),s => s(5)(31),lamdaOut => P(4)(63));
U_F564: entity F port map(lamdaA => P(5)(64),lamdaB => P(5)(96),lamdaOut => P(4)(64));
U_F565: entity F port map(lamdaA => P(5)(65),lamdaB => P(5)(97),lamdaOut => P(4)(65));
U_F566: entity F port map(lamdaA => P(5)(66),lamdaB => P(5)(98),lamdaOut => P(4)(66));
U_F567: entity F port map(lamdaA => P(5)(67),lamdaB => P(5)(99),lamdaOut => P(4)(67));
U_F568: entity F port map(lamdaA => P(5)(68),lamdaB => P(5)(100),lamdaOut => P(4)(68));
U_F569: entity F port map(lamdaA => P(5)(69),lamdaB => P(5)(101),lamdaOut => P(4)(69));
U_F570: entity F port map(lamdaA => P(5)(70),lamdaB => P(5)(102),lamdaOut => P(4)(70));
U_F571: entity F port map(lamdaA => P(5)(71),lamdaB => P(5)(103),lamdaOut => P(4)(71));
U_F572: entity F port map(lamdaA => P(5)(72),lamdaB => P(5)(104),lamdaOut => P(4)(72));
U_F573: entity F port map(lamdaA => P(5)(73),lamdaB => P(5)(105),lamdaOut => P(4)(73));
U_F574: entity F port map(lamdaA => P(5)(74),lamdaB => P(5)(106),lamdaOut => P(4)(74));
U_F575: entity F port map(lamdaA => P(5)(75),lamdaB => P(5)(107),lamdaOut => P(4)(75));
U_F576: entity F port map(lamdaA => P(5)(76),lamdaB => P(5)(108),lamdaOut => P(4)(76));
U_F577: entity F port map(lamdaA => P(5)(77),lamdaB => P(5)(109),lamdaOut => P(4)(77));
U_F578: entity F port map(lamdaA => P(5)(78),lamdaB => P(5)(110),lamdaOut => P(4)(78));
U_F579: entity F port map(lamdaA => P(5)(79),lamdaB => P(5)(111),lamdaOut => P(4)(79));
U_F580: entity F port map(lamdaA => P(5)(80),lamdaB => P(5)(112),lamdaOut => P(4)(80));
U_F581: entity F port map(lamdaA => P(5)(81),lamdaB => P(5)(113),lamdaOut => P(4)(81));
U_F582: entity F port map(lamdaA => P(5)(82),lamdaB => P(5)(114),lamdaOut => P(4)(82));
U_F583: entity F port map(lamdaA => P(5)(83),lamdaB => P(5)(115),lamdaOut => P(4)(83));
U_F584: entity F port map(lamdaA => P(5)(84),lamdaB => P(5)(116),lamdaOut => P(4)(84));
U_F585: entity F port map(lamdaA => P(5)(85),lamdaB => P(5)(117),lamdaOut => P(4)(85));
U_F586: entity F port map(lamdaA => P(5)(86),lamdaB => P(5)(118),lamdaOut => P(4)(86));
U_F587: entity F port map(lamdaA => P(5)(87),lamdaB => P(5)(119),lamdaOut => P(4)(87));
U_F588: entity F port map(lamdaA => P(5)(88),lamdaB => P(5)(120),lamdaOut => P(4)(88));
U_F589: entity F port map(lamdaA => P(5)(89),lamdaB => P(5)(121),lamdaOut => P(4)(89));
U_F590: entity F port map(lamdaA => P(5)(90),lamdaB => P(5)(122),lamdaOut => P(4)(90));
U_F591: entity F port map(lamdaA => P(5)(91),lamdaB => P(5)(123),lamdaOut => P(4)(91));
U_F592: entity F port map(lamdaA => P(5)(92),lamdaB => P(5)(124),lamdaOut => P(4)(92));
U_F593: entity F port map(lamdaA => P(5)(93),lamdaB => P(5)(125),lamdaOut => P(4)(93));
U_F594: entity F port map(lamdaA => P(5)(94),lamdaB => P(5)(126),lamdaOut => P(4)(94));
U_F595: entity F port map(lamdaA => P(5)(95),lamdaB => P(5)(127),lamdaOut => P(4)(95));
U_G596: entity G port map(lamdaA => P(5)(64),lamdaB => P(5)(96),s => s(5)(32),lamdaOut => P(4)(96));
U_G597: entity G port map(lamdaA => P(5)(65),lamdaB => P(5)(97),s => s(5)(33),lamdaOut => P(4)(97));
U_G598: entity G port map(lamdaA => P(5)(66),lamdaB => P(5)(98),s => s(5)(34),lamdaOut => P(4)(98));
U_G599: entity G port map(lamdaA => P(5)(67),lamdaB => P(5)(99),s => s(5)(35),lamdaOut => P(4)(99));
U_G5100: entity G port map(lamdaA => P(5)(68),lamdaB => P(5)(100),s => s(5)(36),lamdaOut => P(4)(100));
U_G5101: entity G port map(lamdaA => P(5)(69),lamdaB => P(5)(101),s => s(5)(37),lamdaOut => P(4)(101));
U_G5102: entity G port map(lamdaA => P(5)(70),lamdaB => P(5)(102),s => s(5)(38),lamdaOut => P(4)(102));
U_G5103: entity G port map(lamdaA => P(5)(71),lamdaB => P(5)(103),s => s(5)(39),lamdaOut => P(4)(103));
U_G5104: entity G port map(lamdaA => P(5)(72),lamdaB => P(5)(104),s => s(5)(40),lamdaOut => P(4)(104));
U_G5105: entity G port map(lamdaA => P(5)(73),lamdaB => P(5)(105),s => s(5)(41),lamdaOut => P(4)(105));
U_G5106: entity G port map(lamdaA => P(5)(74),lamdaB => P(5)(106),s => s(5)(42),lamdaOut => P(4)(106));
U_G5107: entity G port map(lamdaA => P(5)(75),lamdaB => P(5)(107),s => s(5)(43),lamdaOut => P(4)(107));
U_G5108: entity G port map(lamdaA => P(5)(76),lamdaB => P(5)(108),s => s(5)(44),lamdaOut => P(4)(108));
U_G5109: entity G port map(lamdaA => P(5)(77),lamdaB => P(5)(109),s => s(5)(45),lamdaOut => P(4)(109));
U_G5110: entity G port map(lamdaA => P(5)(78),lamdaB => P(5)(110),s => s(5)(46),lamdaOut => P(4)(110));
U_G5111: entity G port map(lamdaA => P(5)(79),lamdaB => P(5)(111),s => s(5)(47),lamdaOut => P(4)(111));
U_G5112: entity G port map(lamdaA => P(5)(80),lamdaB => P(5)(112),s => s(5)(48),lamdaOut => P(4)(112));
U_G5113: entity G port map(lamdaA => P(5)(81),lamdaB => P(5)(113),s => s(5)(49),lamdaOut => P(4)(113));
U_G5114: entity G port map(lamdaA => P(5)(82),lamdaB => P(5)(114),s => s(5)(50),lamdaOut => P(4)(114));
U_G5115: entity G port map(lamdaA => P(5)(83),lamdaB => P(5)(115),s => s(5)(51),lamdaOut => P(4)(115));
U_G5116: entity G port map(lamdaA => P(5)(84),lamdaB => P(5)(116),s => s(5)(52),lamdaOut => P(4)(116));
U_G5117: entity G port map(lamdaA => P(5)(85),lamdaB => P(5)(117),s => s(5)(53),lamdaOut => P(4)(117));
U_G5118: entity G port map(lamdaA => P(5)(86),lamdaB => P(5)(118),s => s(5)(54),lamdaOut => P(4)(118));
U_G5119: entity G port map(lamdaA => P(5)(87),lamdaB => P(5)(119),s => s(5)(55),lamdaOut => P(4)(119));
U_G5120: entity G port map(lamdaA => P(5)(88),lamdaB => P(5)(120),s => s(5)(56),lamdaOut => P(4)(120));
U_G5121: entity G port map(lamdaA => P(5)(89),lamdaB => P(5)(121),s => s(5)(57),lamdaOut => P(4)(121));
U_G5122: entity G port map(lamdaA => P(5)(90),lamdaB => P(5)(122),s => s(5)(58),lamdaOut => P(4)(122));
U_G5123: entity G port map(lamdaA => P(5)(91),lamdaB => P(5)(123),s => s(5)(59),lamdaOut => P(4)(123));
U_G5124: entity G port map(lamdaA => P(5)(92),lamdaB => P(5)(124),s => s(5)(60),lamdaOut => P(4)(124));
U_G5125: entity G port map(lamdaA => P(5)(93),lamdaB => P(5)(125),s => s(5)(61),lamdaOut => P(4)(125));
U_G5126: entity G port map(lamdaA => P(5)(94),lamdaB => P(5)(126),s => s(5)(62),lamdaOut => P(4)(126));
U_G5127: entity G port map(lamdaA => P(5)(95),lamdaB => P(5)(127),s => s(5)(63),lamdaOut => P(4)(127));
U_F5128: entity F port map(lamdaA => P(5)(128),lamdaB => P(5)(160),lamdaOut => P(4)(128));
U_F5129: entity F port map(lamdaA => P(5)(129),lamdaB => P(5)(161),lamdaOut => P(4)(129));
U_F5130: entity F port map(lamdaA => P(5)(130),lamdaB => P(5)(162),lamdaOut => P(4)(130));
U_F5131: entity F port map(lamdaA => P(5)(131),lamdaB => P(5)(163),lamdaOut => P(4)(131));
U_F5132: entity F port map(lamdaA => P(5)(132),lamdaB => P(5)(164),lamdaOut => P(4)(132));
U_F5133: entity F port map(lamdaA => P(5)(133),lamdaB => P(5)(165),lamdaOut => P(4)(133));
U_F5134: entity F port map(lamdaA => P(5)(134),lamdaB => P(5)(166),lamdaOut => P(4)(134));
U_F5135: entity F port map(lamdaA => P(5)(135),lamdaB => P(5)(167),lamdaOut => P(4)(135));
U_F5136: entity F port map(lamdaA => P(5)(136),lamdaB => P(5)(168),lamdaOut => P(4)(136));
U_F5137: entity F port map(lamdaA => P(5)(137),lamdaB => P(5)(169),lamdaOut => P(4)(137));
U_F5138: entity F port map(lamdaA => P(5)(138),lamdaB => P(5)(170),lamdaOut => P(4)(138));
U_F5139: entity F port map(lamdaA => P(5)(139),lamdaB => P(5)(171),lamdaOut => P(4)(139));
U_F5140: entity F port map(lamdaA => P(5)(140),lamdaB => P(5)(172),lamdaOut => P(4)(140));
U_F5141: entity F port map(lamdaA => P(5)(141),lamdaB => P(5)(173),lamdaOut => P(4)(141));
U_F5142: entity F port map(lamdaA => P(5)(142),lamdaB => P(5)(174),lamdaOut => P(4)(142));
U_F5143: entity F port map(lamdaA => P(5)(143),lamdaB => P(5)(175),lamdaOut => P(4)(143));
U_F5144: entity F port map(lamdaA => P(5)(144),lamdaB => P(5)(176),lamdaOut => P(4)(144));
U_F5145: entity F port map(lamdaA => P(5)(145),lamdaB => P(5)(177),lamdaOut => P(4)(145));
U_F5146: entity F port map(lamdaA => P(5)(146),lamdaB => P(5)(178),lamdaOut => P(4)(146));
U_F5147: entity F port map(lamdaA => P(5)(147),lamdaB => P(5)(179),lamdaOut => P(4)(147));
U_F5148: entity F port map(lamdaA => P(5)(148),lamdaB => P(5)(180),lamdaOut => P(4)(148));
U_F5149: entity F port map(lamdaA => P(5)(149),lamdaB => P(5)(181),lamdaOut => P(4)(149));
U_F5150: entity F port map(lamdaA => P(5)(150),lamdaB => P(5)(182),lamdaOut => P(4)(150));
U_F5151: entity F port map(lamdaA => P(5)(151),lamdaB => P(5)(183),lamdaOut => P(4)(151));
U_F5152: entity F port map(lamdaA => P(5)(152),lamdaB => P(5)(184),lamdaOut => P(4)(152));
U_F5153: entity F port map(lamdaA => P(5)(153),lamdaB => P(5)(185),lamdaOut => P(4)(153));
U_F5154: entity F port map(lamdaA => P(5)(154),lamdaB => P(5)(186),lamdaOut => P(4)(154));
U_F5155: entity F port map(lamdaA => P(5)(155),lamdaB => P(5)(187),lamdaOut => P(4)(155));
U_F5156: entity F port map(lamdaA => P(5)(156),lamdaB => P(5)(188),lamdaOut => P(4)(156));
U_F5157: entity F port map(lamdaA => P(5)(157),lamdaB => P(5)(189),lamdaOut => P(4)(157));
U_F5158: entity F port map(lamdaA => P(5)(158),lamdaB => P(5)(190),lamdaOut => P(4)(158));
U_F5159: entity F port map(lamdaA => P(5)(159),lamdaB => P(5)(191),lamdaOut => P(4)(159));
U_G5160: entity G port map(lamdaA => P(5)(128),lamdaB => P(5)(160),s => s(5)(64),lamdaOut => P(4)(160));
U_G5161: entity G port map(lamdaA => P(5)(129),lamdaB => P(5)(161),s => s(5)(65),lamdaOut => P(4)(161));
U_G5162: entity G port map(lamdaA => P(5)(130),lamdaB => P(5)(162),s => s(5)(66),lamdaOut => P(4)(162));
U_G5163: entity G port map(lamdaA => P(5)(131),lamdaB => P(5)(163),s => s(5)(67),lamdaOut => P(4)(163));
U_G5164: entity G port map(lamdaA => P(5)(132),lamdaB => P(5)(164),s => s(5)(68),lamdaOut => P(4)(164));
U_G5165: entity G port map(lamdaA => P(5)(133),lamdaB => P(5)(165),s => s(5)(69),lamdaOut => P(4)(165));
U_G5166: entity G port map(lamdaA => P(5)(134),lamdaB => P(5)(166),s => s(5)(70),lamdaOut => P(4)(166));
U_G5167: entity G port map(lamdaA => P(5)(135),lamdaB => P(5)(167),s => s(5)(71),lamdaOut => P(4)(167));
U_G5168: entity G port map(lamdaA => P(5)(136),lamdaB => P(5)(168),s => s(5)(72),lamdaOut => P(4)(168));
U_G5169: entity G port map(lamdaA => P(5)(137),lamdaB => P(5)(169),s => s(5)(73),lamdaOut => P(4)(169));
U_G5170: entity G port map(lamdaA => P(5)(138),lamdaB => P(5)(170),s => s(5)(74),lamdaOut => P(4)(170));
U_G5171: entity G port map(lamdaA => P(5)(139),lamdaB => P(5)(171),s => s(5)(75),lamdaOut => P(4)(171));
U_G5172: entity G port map(lamdaA => P(5)(140),lamdaB => P(5)(172),s => s(5)(76),lamdaOut => P(4)(172));
U_G5173: entity G port map(lamdaA => P(5)(141),lamdaB => P(5)(173),s => s(5)(77),lamdaOut => P(4)(173));
U_G5174: entity G port map(lamdaA => P(5)(142),lamdaB => P(5)(174),s => s(5)(78),lamdaOut => P(4)(174));
U_G5175: entity G port map(lamdaA => P(5)(143),lamdaB => P(5)(175),s => s(5)(79),lamdaOut => P(4)(175));
U_G5176: entity G port map(lamdaA => P(5)(144),lamdaB => P(5)(176),s => s(5)(80),lamdaOut => P(4)(176));
U_G5177: entity G port map(lamdaA => P(5)(145),lamdaB => P(5)(177),s => s(5)(81),lamdaOut => P(4)(177));
U_G5178: entity G port map(lamdaA => P(5)(146),lamdaB => P(5)(178),s => s(5)(82),lamdaOut => P(4)(178));
U_G5179: entity G port map(lamdaA => P(5)(147),lamdaB => P(5)(179),s => s(5)(83),lamdaOut => P(4)(179));
U_G5180: entity G port map(lamdaA => P(5)(148),lamdaB => P(5)(180),s => s(5)(84),lamdaOut => P(4)(180));
U_G5181: entity G port map(lamdaA => P(5)(149),lamdaB => P(5)(181),s => s(5)(85),lamdaOut => P(4)(181));
U_G5182: entity G port map(lamdaA => P(5)(150),lamdaB => P(5)(182),s => s(5)(86),lamdaOut => P(4)(182));
U_G5183: entity G port map(lamdaA => P(5)(151),lamdaB => P(5)(183),s => s(5)(87),lamdaOut => P(4)(183));
U_G5184: entity G port map(lamdaA => P(5)(152),lamdaB => P(5)(184),s => s(5)(88),lamdaOut => P(4)(184));
U_G5185: entity G port map(lamdaA => P(5)(153),lamdaB => P(5)(185),s => s(5)(89),lamdaOut => P(4)(185));
U_G5186: entity G port map(lamdaA => P(5)(154),lamdaB => P(5)(186),s => s(5)(90),lamdaOut => P(4)(186));
U_G5187: entity G port map(lamdaA => P(5)(155),lamdaB => P(5)(187),s => s(5)(91),lamdaOut => P(4)(187));
U_G5188: entity G port map(lamdaA => P(5)(156),lamdaB => P(5)(188),s => s(5)(92),lamdaOut => P(4)(188));
U_G5189: entity G port map(lamdaA => P(5)(157),lamdaB => P(5)(189),s => s(5)(93),lamdaOut => P(4)(189));
U_G5190: entity G port map(lamdaA => P(5)(158),lamdaB => P(5)(190),s => s(5)(94),lamdaOut => P(4)(190));
U_G5191: entity G port map(lamdaA => P(5)(159),lamdaB => P(5)(191),s => s(5)(95),lamdaOut => P(4)(191));
U_F5192: entity F port map(lamdaA => P(5)(192),lamdaB => P(5)(224),lamdaOut => P(4)(192));
U_F5193: entity F port map(lamdaA => P(5)(193),lamdaB => P(5)(225),lamdaOut => P(4)(193));
U_F5194: entity F port map(lamdaA => P(5)(194),lamdaB => P(5)(226),lamdaOut => P(4)(194));
U_F5195: entity F port map(lamdaA => P(5)(195),lamdaB => P(5)(227),lamdaOut => P(4)(195));
U_F5196: entity F port map(lamdaA => P(5)(196),lamdaB => P(5)(228),lamdaOut => P(4)(196));
U_F5197: entity F port map(lamdaA => P(5)(197),lamdaB => P(5)(229),lamdaOut => P(4)(197));
U_F5198: entity F port map(lamdaA => P(5)(198),lamdaB => P(5)(230),lamdaOut => P(4)(198));
U_F5199: entity F port map(lamdaA => P(5)(199),lamdaB => P(5)(231),lamdaOut => P(4)(199));
U_F5200: entity F port map(lamdaA => P(5)(200),lamdaB => P(5)(232),lamdaOut => P(4)(200));
U_F5201: entity F port map(lamdaA => P(5)(201),lamdaB => P(5)(233),lamdaOut => P(4)(201));
U_F5202: entity F port map(lamdaA => P(5)(202),lamdaB => P(5)(234),lamdaOut => P(4)(202));
U_F5203: entity F port map(lamdaA => P(5)(203),lamdaB => P(5)(235),lamdaOut => P(4)(203));
U_F5204: entity F port map(lamdaA => P(5)(204),lamdaB => P(5)(236),lamdaOut => P(4)(204));
U_F5205: entity F port map(lamdaA => P(5)(205),lamdaB => P(5)(237),lamdaOut => P(4)(205));
U_F5206: entity F port map(lamdaA => P(5)(206),lamdaB => P(5)(238),lamdaOut => P(4)(206));
U_F5207: entity F port map(lamdaA => P(5)(207),lamdaB => P(5)(239),lamdaOut => P(4)(207));
U_F5208: entity F port map(lamdaA => P(5)(208),lamdaB => P(5)(240),lamdaOut => P(4)(208));
U_F5209: entity F port map(lamdaA => P(5)(209),lamdaB => P(5)(241),lamdaOut => P(4)(209));
U_F5210: entity F port map(lamdaA => P(5)(210),lamdaB => P(5)(242),lamdaOut => P(4)(210));
U_F5211: entity F port map(lamdaA => P(5)(211),lamdaB => P(5)(243),lamdaOut => P(4)(211));
U_F5212: entity F port map(lamdaA => P(5)(212),lamdaB => P(5)(244),lamdaOut => P(4)(212));
U_F5213: entity F port map(lamdaA => P(5)(213),lamdaB => P(5)(245),lamdaOut => P(4)(213));
U_F5214: entity F port map(lamdaA => P(5)(214),lamdaB => P(5)(246),lamdaOut => P(4)(214));
U_F5215: entity F port map(lamdaA => P(5)(215),lamdaB => P(5)(247),lamdaOut => P(4)(215));
U_F5216: entity F port map(lamdaA => P(5)(216),lamdaB => P(5)(248),lamdaOut => P(4)(216));
U_F5217: entity F port map(lamdaA => P(5)(217),lamdaB => P(5)(249),lamdaOut => P(4)(217));
U_F5218: entity F port map(lamdaA => P(5)(218),lamdaB => P(5)(250),lamdaOut => P(4)(218));
U_F5219: entity F port map(lamdaA => P(5)(219),lamdaB => P(5)(251),lamdaOut => P(4)(219));
U_F5220: entity F port map(lamdaA => P(5)(220),lamdaB => P(5)(252),lamdaOut => P(4)(220));
U_F5221: entity F port map(lamdaA => P(5)(221),lamdaB => P(5)(253),lamdaOut => P(4)(221));
U_F5222: entity F port map(lamdaA => P(5)(222),lamdaB => P(5)(254),lamdaOut => P(4)(222));
U_F5223: entity F port map(lamdaA => P(5)(223),lamdaB => P(5)(255),lamdaOut => P(4)(223));
U_G5224: entity G port map(lamdaA => P(5)(192),lamdaB => P(5)(224),s => s(5)(96),lamdaOut => P(4)(224));
U_G5225: entity G port map(lamdaA => P(5)(193),lamdaB => P(5)(225),s => s(5)(97),lamdaOut => P(4)(225));
U_G5226: entity G port map(lamdaA => P(5)(194),lamdaB => P(5)(226),s => s(5)(98),lamdaOut => P(4)(226));
U_G5227: entity G port map(lamdaA => P(5)(195),lamdaB => P(5)(227),s => s(5)(99),lamdaOut => P(4)(227));
U_G5228: entity G port map(lamdaA => P(5)(196),lamdaB => P(5)(228),s => s(5)(100),lamdaOut => P(4)(228));
U_G5229: entity G port map(lamdaA => P(5)(197),lamdaB => P(5)(229),s => s(5)(101),lamdaOut => P(4)(229));
U_G5230: entity G port map(lamdaA => P(5)(198),lamdaB => P(5)(230),s => s(5)(102),lamdaOut => P(4)(230));
U_G5231: entity G port map(lamdaA => P(5)(199),lamdaB => P(5)(231),s => s(5)(103),lamdaOut => P(4)(231));
U_G5232: entity G port map(lamdaA => P(5)(200),lamdaB => P(5)(232),s => s(5)(104),lamdaOut => P(4)(232));
U_G5233: entity G port map(lamdaA => P(5)(201),lamdaB => P(5)(233),s => s(5)(105),lamdaOut => P(4)(233));
U_G5234: entity G port map(lamdaA => P(5)(202),lamdaB => P(5)(234),s => s(5)(106),lamdaOut => P(4)(234));
U_G5235: entity G port map(lamdaA => P(5)(203),lamdaB => P(5)(235),s => s(5)(107),lamdaOut => P(4)(235));
U_G5236: entity G port map(lamdaA => P(5)(204),lamdaB => P(5)(236),s => s(5)(108),lamdaOut => P(4)(236));
U_G5237: entity G port map(lamdaA => P(5)(205),lamdaB => P(5)(237),s => s(5)(109),lamdaOut => P(4)(237));
U_G5238: entity G port map(lamdaA => P(5)(206),lamdaB => P(5)(238),s => s(5)(110),lamdaOut => P(4)(238));
U_G5239: entity G port map(lamdaA => P(5)(207),lamdaB => P(5)(239),s => s(5)(111),lamdaOut => P(4)(239));
U_G5240: entity G port map(lamdaA => P(5)(208),lamdaB => P(5)(240),s => s(5)(112),lamdaOut => P(4)(240));
U_G5241: entity G port map(lamdaA => P(5)(209),lamdaB => P(5)(241),s => s(5)(113),lamdaOut => P(4)(241));
U_G5242: entity G port map(lamdaA => P(5)(210),lamdaB => P(5)(242),s => s(5)(114),lamdaOut => P(4)(242));
U_G5243: entity G port map(lamdaA => P(5)(211),lamdaB => P(5)(243),s => s(5)(115),lamdaOut => P(4)(243));
U_G5244: entity G port map(lamdaA => P(5)(212),lamdaB => P(5)(244),s => s(5)(116),lamdaOut => P(4)(244));
U_G5245: entity G port map(lamdaA => P(5)(213),lamdaB => P(5)(245),s => s(5)(117),lamdaOut => P(4)(245));
U_G5246: entity G port map(lamdaA => P(5)(214),lamdaB => P(5)(246),s => s(5)(118),lamdaOut => P(4)(246));
U_G5247: entity G port map(lamdaA => P(5)(215),lamdaB => P(5)(247),s => s(5)(119),lamdaOut => P(4)(247));
U_G5248: entity G port map(lamdaA => P(5)(216),lamdaB => P(5)(248),s => s(5)(120),lamdaOut => P(4)(248));
U_G5249: entity G port map(lamdaA => P(5)(217),lamdaB => P(5)(249),s => s(5)(121),lamdaOut => P(4)(249));
U_G5250: entity G port map(lamdaA => P(5)(218),lamdaB => P(5)(250),s => s(5)(122),lamdaOut => P(4)(250));
U_G5251: entity G port map(lamdaA => P(5)(219),lamdaB => P(5)(251),s => s(5)(123),lamdaOut => P(4)(251));
U_G5252: entity G port map(lamdaA => P(5)(220),lamdaB => P(5)(252),s => s(5)(124),lamdaOut => P(4)(252));
U_G5253: entity G port map(lamdaA => P(5)(221),lamdaB => P(5)(253),s => s(5)(125),lamdaOut => P(4)(253));
U_G5254: entity G port map(lamdaA => P(5)(222),lamdaB => P(5)(254),s => s(5)(126),lamdaOut => P(4)(254));
U_G5255: entity G port map(lamdaA => P(5)(223),lamdaB => P(5)(255),s => s(5)(127),lamdaOut => P(4)(255));
U_F5256: entity F port map(lamdaA => P(5)(256),lamdaB => P(5)(288),lamdaOut => P(4)(256));
U_F5257: entity F port map(lamdaA => P(5)(257),lamdaB => P(5)(289),lamdaOut => P(4)(257));
U_F5258: entity F port map(lamdaA => P(5)(258),lamdaB => P(5)(290),lamdaOut => P(4)(258));
U_F5259: entity F port map(lamdaA => P(5)(259),lamdaB => P(5)(291),lamdaOut => P(4)(259));
U_F5260: entity F port map(lamdaA => P(5)(260),lamdaB => P(5)(292),lamdaOut => P(4)(260));
U_F5261: entity F port map(lamdaA => P(5)(261),lamdaB => P(5)(293),lamdaOut => P(4)(261));
U_F5262: entity F port map(lamdaA => P(5)(262),lamdaB => P(5)(294),lamdaOut => P(4)(262));
U_F5263: entity F port map(lamdaA => P(5)(263),lamdaB => P(5)(295),lamdaOut => P(4)(263));
U_F5264: entity F port map(lamdaA => P(5)(264),lamdaB => P(5)(296),lamdaOut => P(4)(264));
U_F5265: entity F port map(lamdaA => P(5)(265),lamdaB => P(5)(297),lamdaOut => P(4)(265));
U_F5266: entity F port map(lamdaA => P(5)(266),lamdaB => P(5)(298),lamdaOut => P(4)(266));
U_F5267: entity F port map(lamdaA => P(5)(267),lamdaB => P(5)(299),lamdaOut => P(4)(267));
U_F5268: entity F port map(lamdaA => P(5)(268),lamdaB => P(5)(300),lamdaOut => P(4)(268));
U_F5269: entity F port map(lamdaA => P(5)(269),lamdaB => P(5)(301),lamdaOut => P(4)(269));
U_F5270: entity F port map(lamdaA => P(5)(270),lamdaB => P(5)(302),lamdaOut => P(4)(270));
U_F5271: entity F port map(lamdaA => P(5)(271),lamdaB => P(5)(303),lamdaOut => P(4)(271));
U_F5272: entity F port map(lamdaA => P(5)(272),lamdaB => P(5)(304),lamdaOut => P(4)(272));
U_F5273: entity F port map(lamdaA => P(5)(273),lamdaB => P(5)(305),lamdaOut => P(4)(273));
U_F5274: entity F port map(lamdaA => P(5)(274),lamdaB => P(5)(306),lamdaOut => P(4)(274));
U_F5275: entity F port map(lamdaA => P(5)(275),lamdaB => P(5)(307),lamdaOut => P(4)(275));
U_F5276: entity F port map(lamdaA => P(5)(276),lamdaB => P(5)(308),lamdaOut => P(4)(276));
U_F5277: entity F port map(lamdaA => P(5)(277),lamdaB => P(5)(309),lamdaOut => P(4)(277));
U_F5278: entity F port map(lamdaA => P(5)(278),lamdaB => P(5)(310),lamdaOut => P(4)(278));
U_F5279: entity F port map(lamdaA => P(5)(279),lamdaB => P(5)(311),lamdaOut => P(4)(279));
U_F5280: entity F port map(lamdaA => P(5)(280),lamdaB => P(5)(312),lamdaOut => P(4)(280));
U_F5281: entity F port map(lamdaA => P(5)(281),lamdaB => P(5)(313),lamdaOut => P(4)(281));
U_F5282: entity F port map(lamdaA => P(5)(282),lamdaB => P(5)(314),lamdaOut => P(4)(282));
U_F5283: entity F port map(lamdaA => P(5)(283),lamdaB => P(5)(315),lamdaOut => P(4)(283));
U_F5284: entity F port map(lamdaA => P(5)(284),lamdaB => P(5)(316),lamdaOut => P(4)(284));
U_F5285: entity F port map(lamdaA => P(5)(285),lamdaB => P(5)(317),lamdaOut => P(4)(285));
U_F5286: entity F port map(lamdaA => P(5)(286),lamdaB => P(5)(318),lamdaOut => P(4)(286));
U_F5287: entity F port map(lamdaA => P(5)(287),lamdaB => P(5)(319),lamdaOut => P(4)(287));
U_G5288: entity G port map(lamdaA => P(5)(256),lamdaB => P(5)(288),s => s(5)(128),lamdaOut => P(4)(288));
U_G5289: entity G port map(lamdaA => P(5)(257),lamdaB => P(5)(289),s => s(5)(129),lamdaOut => P(4)(289));
U_G5290: entity G port map(lamdaA => P(5)(258),lamdaB => P(5)(290),s => s(5)(130),lamdaOut => P(4)(290));
U_G5291: entity G port map(lamdaA => P(5)(259),lamdaB => P(5)(291),s => s(5)(131),lamdaOut => P(4)(291));
U_G5292: entity G port map(lamdaA => P(5)(260),lamdaB => P(5)(292),s => s(5)(132),lamdaOut => P(4)(292));
U_G5293: entity G port map(lamdaA => P(5)(261),lamdaB => P(5)(293),s => s(5)(133),lamdaOut => P(4)(293));
U_G5294: entity G port map(lamdaA => P(5)(262),lamdaB => P(5)(294),s => s(5)(134),lamdaOut => P(4)(294));
U_G5295: entity G port map(lamdaA => P(5)(263),lamdaB => P(5)(295),s => s(5)(135),lamdaOut => P(4)(295));
U_G5296: entity G port map(lamdaA => P(5)(264),lamdaB => P(5)(296),s => s(5)(136),lamdaOut => P(4)(296));
U_G5297: entity G port map(lamdaA => P(5)(265),lamdaB => P(5)(297),s => s(5)(137),lamdaOut => P(4)(297));
U_G5298: entity G port map(lamdaA => P(5)(266),lamdaB => P(5)(298),s => s(5)(138),lamdaOut => P(4)(298));
U_G5299: entity G port map(lamdaA => P(5)(267),lamdaB => P(5)(299),s => s(5)(139),lamdaOut => P(4)(299));
U_G5300: entity G port map(lamdaA => P(5)(268),lamdaB => P(5)(300),s => s(5)(140),lamdaOut => P(4)(300));
U_G5301: entity G port map(lamdaA => P(5)(269),lamdaB => P(5)(301),s => s(5)(141),lamdaOut => P(4)(301));
U_G5302: entity G port map(lamdaA => P(5)(270),lamdaB => P(5)(302),s => s(5)(142),lamdaOut => P(4)(302));
U_G5303: entity G port map(lamdaA => P(5)(271),lamdaB => P(5)(303),s => s(5)(143),lamdaOut => P(4)(303));
U_G5304: entity G port map(lamdaA => P(5)(272),lamdaB => P(5)(304),s => s(5)(144),lamdaOut => P(4)(304));
U_G5305: entity G port map(lamdaA => P(5)(273),lamdaB => P(5)(305),s => s(5)(145),lamdaOut => P(4)(305));
U_G5306: entity G port map(lamdaA => P(5)(274),lamdaB => P(5)(306),s => s(5)(146),lamdaOut => P(4)(306));
U_G5307: entity G port map(lamdaA => P(5)(275),lamdaB => P(5)(307),s => s(5)(147),lamdaOut => P(4)(307));
U_G5308: entity G port map(lamdaA => P(5)(276),lamdaB => P(5)(308),s => s(5)(148),lamdaOut => P(4)(308));
U_G5309: entity G port map(lamdaA => P(5)(277),lamdaB => P(5)(309),s => s(5)(149),lamdaOut => P(4)(309));
U_G5310: entity G port map(lamdaA => P(5)(278),lamdaB => P(5)(310),s => s(5)(150),lamdaOut => P(4)(310));
U_G5311: entity G port map(lamdaA => P(5)(279),lamdaB => P(5)(311),s => s(5)(151),lamdaOut => P(4)(311));
U_G5312: entity G port map(lamdaA => P(5)(280),lamdaB => P(5)(312),s => s(5)(152),lamdaOut => P(4)(312));
U_G5313: entity G port map(lamdaA => P(5)(281),lamdaB => P(5)(313),s => s(5)(153),lamdaOut => P(4)(313));
U_G5314: entity G port map(lamdaA => P(5)(282),lamdaB => P(5)(314),s => s(5)(154),lamdaOut => P(4)(314));
U_G5315: entity G port map(lamdaA => P(5)(283),lamdaB => P(5)(315),s => s(5)(155),lamdaOut => P(4)(315));
U_G5316: entity G port map(lamdaA => P(5)(284),lamdaB => P(5)(316),s => s(5)(156),lamdaOut => P(4)(316));
U_G5317: entity G port map(lamdaA => P(5)(285),lamdaB => P(5)(317),s => s(5)(157),lamdaOut => P(4)(317));
U_G5318: entity G port map(lamdaA => P(5)(286),lamdaB => P(5)(318),s => s(5)(158),lamdaOut => P(4)(318));
U_G5319: entity G port map(lamdaA => P(5)(287),lamdaB => P(5)(319),s => s(5)(159),lamdaOut => P(4)(319));
U_F5320: entity F port map(lamdaA => P(5)(320),lamdaB => P(5)(352),lamdaOut => P(4)(320));
U_F5321: entity F port map(lamdaA => P(5)(321),lamdaB => P(5)(353),lamdaOut => P(4)(321));
U_F5322: entity F port map(lamdaA => P(5)(322),lamdaB => P(5)(354),lamdaOut => P(4)(322));
U_F5323: entity F port map(lamdaA => P(5)(323),lamdaB => P(5)(355),lamdaOut => P(4)(323));
U_F5324: entity F port map(lamdaA => P(5)(324),lamdaB => P(5)(356),lamdaOut => P(4)(324));
U_F5325: entity F port map(lamdaA => P(5)(325),lamdaB => P(5)(357),lamdaOut => P(4)(325));
U_F5326: entity F port map(lamdaA => P(5)(326),lamdaB => P(5)(358),lamdaOut => P(4)(326));
U_F5327: entity F port map(lamdaA => P(5)(327),lamdaB => P(5)(359),lamdaOut => P(4)(327));
U_F5328: entity F port map(lamdaA => P(5)(328),lamdaB => P(5)(360),lamdaOut => P(4)(328));
U_F5329: entity F port map(lamdaA => P(5)(329),lamdaB => P(5)(361),lamdaOut => P(4)(329));
U_F5330: entity F port map(lamdaA => P(5)(330),lamdaB => P(5)(362),lamdaOut => P(4)(330));
U_F5331: entity F port map(lamdaA => P(5)(331),lamdaB => P(5)(363),lamdaOut => P(4)(331));
U_F5332: entity F port map(lamdaA => P(5)(332),lamdaB => P(5)(364),lamdaOut => P(4)(332));
U_F5333: entity F port map(lamdaA => P(5)(333),lamdaB => P(5)(365),lamdaOut => P(4)(333));
U_F5334: entity F port map(lamdaA => P(5)(334),lamdaB => P(5)(366),lamdaOut => P(4)(334));
U_F5335: entity F port map(lamdaA => P(5)(335),lamdaB => P(5)(367),lamdaOut => P(4)(335));
U_F5336: entity F port map(lamdaA => P(5)(336),lamdaB => P(5)(368),lamdaOut => P(4)(336));
U_F5337: entity F port map(lamdaA => P(5)(337),lamdaB => P(5)(369),lamdaOut => P(4)(337));
U_F5338: entity F port map(lamdaA => P(5)(338),lamdaB => P(5)(370),lamdaOut => P(4)(338));
U_F5339: entity F port map(lamdaA => P(5)(339),lamdaB => P(5)(371),lamdaOut => P(4)(339));
U_F5340: entity F port map(lamdaA => P(5)(340),lamdaB => P(5)(372),lamdaOut => P(4)(340));
U_F5341: entity F port map(lamdaA => P(5)(341),lamdaB => P(5)(373),lamdaOut => P(4)(341));
U_F5342: entity F port map(lamdaA => P(5)(342),lamdaB => P(5)(374),lamdaOut => P(4)(342));
U_F5343: entity F port map(lamdaA => P(5)(343),lamdaB => P(5)(375),lamdaOut => P(4)(343));
U_F5344: entity F port map(lamdaA => P(5)(344),lamdaB => P(5)(376),lamdaOut => P(4)(344));
U_F5345: entity F port map(lamdaA => P(5)(345),lamdaB => P(5)(377),lamdaOut => P(4)(345));
U_F5346: entity F port map(lamdaA => P(5)(346),lamdaB => P(5)(378),lamdaOut => P(4)(346));
U_F5347: entity F port map(lamdaA => P(5)(347),lamdaB => P(5)(379),lamdaOut => P(4)(347));
U_F5348: entity F port map(lamdaA => P(5)(348),lamdaB => P(5)(380),lamdaOut => P(4)(348));
U_F5349: entity F port map(lamdaA => P(5)(349),lamdaB => P(5)(381),lamdaOut => P(4)(349));
U_F5350: entity F port map(lamdaA => P(5)(350),lamdaB => P(5)(382),lamdaOut => P(4)(350));
U_F5351: entity F port map(lamdaA => P(5)(351),lamdaB => P(5)(383),lamdaOut => P(4)(351));
U_G5352: entity G port map(lamdaA => P(5)(320),lamdaB => P(5)(352),s => s(5)(160),lamdaOut => P(4)(352));
U_G5353: entity G port map(lamdaA => P(5)(321),lamdaB => P(5)(353),s => s(5)(161),lamdaOut => P(4)(353));
U_G5354: entity G port map(lamdaA => P(5)(322),lamdaB => P(5)(354),s => s(5)(162),lamdaOut => P(4)(354));
U_G5355: entity G port map(lamdaA => P(5)(323),lamdaB => P(5)(355),s => s(5)(163),lamdaOut => P(4)(355));
U_G5356: entity G port map(lamdaA => P(5)(324),lamdaB => P(5)(356),s => s(5)(164),lamdaOut => P(4)(356));
U_G5357: entity G port map(lamdaA => P(5)(325),lamdaB => P(5)(357),s => s(5)(165),lamdaOut => P(4)(357));
U_G5358: entity G port map(lamdaA => P(5)(326),lamdaB => P(5)(358),s => s(5)(166),lamdaOut => P(4)(358));
U_G5359: entity G port map(lamdaA => P(5)(327),lamdaB => P(5)(359),s => s(5)(167),lamdaOut => P(4)(359));
U_G5360: entity G port map(lamdaA => P(5)(328),lamdaB => P(5)(360),s => s(5)(168),lamdaOut => P(4)(360));
U_G5361: entity G port map(lamdaA => P(5)(329),lamdaB => P(5)(361),s => s(5)(169),lamdaOut => P(4)(361));
U_G5362: entity G port map(lamdaA => P(5)(330),lamdaB => P(5)(362),s => s(5)(170),lamdaOut => P(4)(362));
U_G5363: entity G port map(lamdaA => P(5)(331),lamdaB => P(5)(363),s => s(5)(171),lamdaOut => P(4)(363));
U_G5364: entity G port map(lamdaA => P(5)(332),lamdaB => P(5)(364),s => s(5)(172),lamdaOut => P(4)(364));
U_G5365: entity G port map(lamdaA => P(5)(333),lamdaB => P(5)(365),s => s(5)(173),lamdaOut => P(4)(365));
U_G5366: entity G port map(lamdaA => P(5)(334),lamdaB => P(5)(366),s => s(5)(174),lamdaOut => P(4)(366));
U_G5367: entity G port map(lamdaA => P(5)(335),lamdaB => P(5)(367),s => s(5)(175),lamdaOut => P(4)(367));
U_G5368: entity G port map(lamdaA => P(5)(336),lamdaB => P(5)(368),s => s(5)(176),lamdaOut => P(4)(368));
U_G5369: entity G port map(lamdaA => P(5)(337),lamdaB => P(5)(369),s => s(5)(177),lamdaOut => P(4)(369));
U_G5370: entity G port map(lamdaA => P(5)(338),lamdaB => P(5)(370),s => s(5)(178),lamdaOut => P(4)(370));
U_G5371: entity G port map(lamdaA => P(5)(339),lamdaB => P(5)(371),s => s(5)(179),lamdaOut => P(4)(371));
U_G5372: entity G port map(lamdaA => P(5)(340),lamdaB => P(5)(372),s => s(5)(180),lamdaOut => P(4)(372));
U_G5373: entity G port map(lamdaA => P(5)(341),lamdaB => P(5)(373),s => s(5)(181),lamdaOut => P(4)(373));
U_G5374: entity G port map(lamdaA => P(5)(342),lamdaB => P(5)(374),s => s(5)(182),lamdaOut => P(4)(374));
U_G5375: entity G port map(lamdaA => P(5)(343),lamdaB => P(5)(375),s => s(5)(183),lamdaOut => P(4)(375));
U_G5376: entity G port map(lamdaA => P(5)(344),lamdaB => P(5)(376),s => s(5)(184),lamdaOut => P(4)(376));
U_G5377: entity G port map(lamdaA => P(5)(345),lamdaB => P(5)(377),s => s(5)(185),lamdaOut => P(4)(377));
U_G5378: entity G port map(lamdaA => P(5)(346),lamdaB => P(5)(378),s => s(5)(186),lamdaOut => P(4)(378));
U_G5379: entity G port map(lamdaA => P(5)(347),lamdaB => P(5)(379),s => s(5)(187),lamdaOut => P(4)(379));
U_G5380: entity G port map(lamdaA => P(5)(348),lamdaB => P(5)(380),s => s(5)(188),lamdaOut => P(4)(380));
U_G5381: entity G port map(lamdaA => P(5)(349),lamdaB => P(5)(381),s => s(5)(189),lamdaOut => P(4)(381));
U_G5382: entity G port map(lamdaA => P(5)(350),lamdaB => P(5)(382),s => s(5)(190),lamdaOut => P(4)(382));
U_G5383: entity G port map(lamdaA => P(5)(351),lamdaB => P(5)(383),s => s(5)(191),lamdaOut => P(4)(383));
U_F5384: entity F port map(lamdaA => P(5)(384),lamdaB => P(5)(416),lamdaOut => P(4)(384));
U_F5385: entity F port map(lamdaA => P(5)(385),lamdaB => P(5)(417),lamdaOut => P(4)(385));
U_F5386: entity F port map(lamdaA => P(5)(386),lamdaB => P(5)(418),lamdaOut => P(4)(386));
U_F5387: entity F port map(lamdaA => P(5)(387),lamdaB => P(5)(419),lamdaOut => P(4)(387));
U_F5388: entity F port map(lamdaA => P(5)(388),lamdaB => P(5)(420),lamdaOut => P(4)(388));
U_F5389: entity F port map(lamdaA => P(5)(389),lamdaB => P(5)(421),lamdaOut => P(4)(389));
U_F5390: entity F port map(lamdaA => P(5)(390),lamdaB => P(5)(422),lamdaOut => P(4)(390));
U_F5391: entity F port map(lamdaA => P(5)(391),lamdaB => P(5)(423),lamdaOut => P(4)(391));
U_F5392: entity F port map(lamdaA => P(5)(392),lamdaB => P(5)(424),lamdaOut => P(4)(392));
U_F5393: entity F port map(lamdaA => P(5)(393),lamdaB => P(5)(425),lamdaOut => P(4)(393));
U_F5394: entity F port map(lamdaA => P(5)(394),lamdaB => P(5)(426),lamdaOut => P(4)(394));
U_F5395: entity F port map(lamdaA => P(5)(395),lamdaB => P(5)(427),lamdaOut => P(4)(395));
U_F5396: entity F port map(lamdaA => P(5)(396),lamdaB => P(5)(428),lamdaOut => P(4)(396));
U_F5397: entity F port map(lamdaA => P(5)(397),lamdaB => P(5)(429),lamdaOut => P(4)(397));
U_F5398: entity F port map(lamdaA => P(5)(398),lamdaB => P(5)(430),lamdaOut => P(4)(398));
U_F5399: entity F port map(lamdaA => P(5)(399),lamdaB => P(5)(431),lamdaOut => P(4)(399));
U_F5400: entity F port map(lamdaA => P(5)(400),lamdaB => P(5)(432),lamdaOut => P(4)(400));
U_F5401: entity F port map(lamdaA => P(5)(401),lamdaB => P(5)(433),lamdaOut => P(4)(401));
U_F5402: entity F port map(lamdaA => P(5)(402),lamdaB => P(5)(434),lamdaOut => P(4)(402));
U_F5403: entity F port map(lamdaA => P(5)(403),lamdaB => P(5)(435),lamdaOut => P(4)(403));
U_F5404: entity F port map(lamdaA => P(5)(404),lamdaB => P(5)(436),lamdaOut => P(4)(404));
U_F5405: entity F port map(lamdaA => P(5)(405),lamdaB => P(5)(437),lamdaOut => P(4)(405));
U_F5406: entity F port map(lamdaA => P(5)(406),lamdaB => P(5)(438),lamdaOut => P(4)(406));
U_F5407: entity F port map(lamdaA => P(5)(407),lamdaB => P(5)(439),lamdaOut => P(4)(407));
U_F5408: entity F port map(lamdaA => P(5)(408),lamdaB => P(5)(440),lamdaOut => P(4)(408));
U_F5409: entity F port map(lamdaA => P(5)(409),lamdaB => P(5)(441),lamdaOut => P(4)(409));
U_F5410: entity F port map(lamdaA => P(5)(410),lamdaB => P(5)(442),lamdaOut => P(4)(410));
U_F5411: entity F port map(lamdaA => P(5)(411),lamdaB => P(5)(443),lamdaOut => P(4)(411));
U_F5412: entity F port map(lamdaA => P(5)(412),lamdaB => P(5)(444),lamdaOut => P(4)(412));
U_F5413: entity F port map(lamdaA => P(5)(413),lamdaB => P(5)(445),lamdaOut => P(4)(413));
U_F5414: entity F port map(lamdaA => P(5)(414),lamdaB => P(5)(446),lamdaOut => P(4)(414));
U_F5415: entity F port map(lamdaA => P(5)(415),lamdaB => P(5)(447),lamdaOut => P(4)(415));
U_G5416: entity G port map(lamdaA => P(5)(384),lamdaB => P(5)(416),s => s(5)(192),lamdaOut => P(4)(416));
U_G5417: entity G port map(lamdaA => P(5)(385),lamdaB => P(5)(417),s => s(5)(193),lamdaOut => P(4)(417));
U_G5418: entity G port map(lamdaA => P(5)(386),lamdaB => P(5)(418),s => s(5)(194),lamdaOut => P(4)(418));
U_G5419: entity G port map(lamdaA => P(5)(387),lamdaB => P(5)(419),s => s(5)(195),lamdaOut => P(4)(419));
U_G5420: entity G port map(lamdaA => P(5)(388),lamdaB => P(5)(420),s => s(5)(196),lamdaOut => P(4)(420));
U_G5421: entity G port map(lamdaA => P(5)(389),lamdaB => P(5)(421),s => s(5)(197),lamdaOut => P(4)(421));
U_G5422: entity G port map(lamdaA => P(5)(390),lamdaB => P(5)(422),s => s(5)(198),lamdaOut => P(4)(422));
U_G5423: entity G port map(lamdaA => P(5)(391),lamdaB => P(5)(423),s => s(5)(199),lamdaOut => P(4)(423));
U_G5424: entity G port map(lamdaA => P(5)(392),lamdaB => P(5)(424),s => s(5)(200),lamdaOut => P(4)(424));
U_G5425: entity G port map(lamdaA => P(5)(393),lamdaB => P(5)(425),s => s(5)(201),lamdaOut => P(4)(425));
U_G5426: entity G port map(lamdaA => P(5)(394),lamdaB => P(5)(426),s => s(5)(202),lamdaOut => P(4)(426));
U_G5427: entity G port map(lamdaA => P(5)(395),lamdaB => P(5)(427),s => s(5)(203),lamdaOut => P(4)(427));
U_G5428: entity G port map(lamdaA => P(5)(396),lamdaB => P(5)(428),s => s(5)(204),lamdaOut => P(4)(428));
U_G5429: entity G port map(lamdaA => P(5)(397),lamdaB => P(5)(429),s => s(5)(205),lamdaOut => P(4)(429));
U_G5430: entity G port map(lamdaA => P(5)(398),lamdaB => P(5)(430),s => s(5)(206),lamdaOut => P(4)(430));
U_G5431: entity G port map(lamdaA => P(5)(399),lamdaB => P(5)(431),s => s(5)(207),lamdaOut => P(4)(431));
U_G5432: entity G port map(lamdaA => P(5)(400),lamdaB => P(5)(432),s => s(5)(208),lamdaOut => P(4)(432));
U_G5433: entity G port map(lamdaA => P(5)(401),lamdaB => P(5)(433),s => s(5)(209),lamdaOut => P(4)(433));
U_G5434: entity G port map(lamdaA => P(5)(402),lamdaB => P(5)(434),s => s(5)(210),lamdaOut => P(4)(434));
U_G5435: entity G port map(lamdaA => P(5)(403),lamdaB => P(5)(435),s => s(5)(211),lamdaOut => P(4)(435));
U_G5436: entity G port map(lamdaA => P(5)(404),lamdaB => P(5)(436),s => s(5)(212),lamdaOut => P(4)(436));
U_G5437: entity G port map(lamdaA => P(5)(405),lamdaB => P(5)(437),s => s(5)(213),lamdaOut => P(4)(437));
U_G5438: entity G port map(lamdaA => P(5)(406),lamdaB => P(5)(438),s => s(5)(214),lamdaOut => P(4)(438));
U_G5439: entity G port map(lamdaA => P(5)(407),lamdaB => P(5)(439),s => s(5)(215),lamdaOut => P(4)(439));
U_G5440: entity G port map(lamdaA => P(5)(408),lamdaB => P(5)(440),s => s(5)(216),lamdaOut => P(4)(440));
U_G5441: entity G port map(lamdaA => P(5)(409),lamdaB => P(5)(441),s => s(5)(217),lamdaOut => P(4)(441));
U_G5442: entity G port map(lamdaA => P(5)(410),lamdaB => P(5)(442),s => s(5)(218),lamdaOut => P(4)(442));
U_G5443: entity G port map(lamdaA => P(5)(411),lamdaB => P(5)(443),s => s(5)(219),lamdaOut => P(4)(443));
U_G5444: entity G port map(lamdaA => P(5)(412),lamdaB => P(5)(444),s => s(5)(220),lamdaOut => P(4)(444));
U_G5445: entity G port map(lamdaA => P(5)(413),lamdaB => P(5)(445),s => s(5)(221),lamdaOut => P(4)(445));
U_G5446: entity G port map(lamdaA => P(5)(414),lamdaB => P(5)(446),s => s(5)(222),lamdaOut => P(4)(446));
U_G5447: entity G port map(lamdaA => P(5)(415),lamdaB => P(5)(447),s => s(5)(223),lamdaOut => P(4)(447));
U_F5448: entity F port map(lamdaA => P(5)(448),lamdaB => P(5)(480),lamdaOut => P(4)(448));
U_F5449: entity F port map(lamdaA => P(5)(449),lamdaB => P(5)(481),lamdaOut => P(4)(449));
U_F5450: entity F port map(lamdaA => P(5)(450),lamdaB => P(5)(482),lamdaOut => P(4)(450));
U_F5451: entity F port map(lamdaA => P(5)(451),lamdaB => P(5)(483),lamdaOut => P(4)(451));
U_F5452: entity F port map(lamdaA => P(5)(452),lamdaB => P(5)(484),lamdaOut => P(4)(452));
U_F5453: entity F port map(lamdaA => P(5)(453),lamdaB => P(5)(485),lamdaOut => P(4)(453));
U_F5454: entity F port map(lamdaA => P(5)(454),lamdaB => P(5)(486),lamdaOut => P(4)(454));
U_F5455: entity F port map(lamdaA => P(5)(455),lamdaB => P(5)(487),lamdaOut => P(4)(455));
U_F5456: entity F port map(lamdaA => P(5)(456),lamdaB => P(5)(488),lamdaOut => P(4)(456));
U_F5457: entity F port map(lamdaA => P(5)(457),lamdaB => P(5)(489),lamdaOut => P(4)(457));
U_F5458: entity F port map(lamdaA => P(5)(458),lamdaB => P(5)(490),lamdaOut => P(4)(458));
U_F5459: entity F port map(lamdaA => P(5)(459),lamdaB => P(5)(491),lamdaOut => P(4)(459));
U_F5460: entity F port map(lamdaA => P(5)(460),lamdaB => P(5)(492),lamdaOut => P(4)(460));
U_F5461: entity F port map(lamdaA => P(5)(461),lamdaB => P(5)(493),lamdaOut => P(4)(461));
U_F5462: entity F port map(lamdaA => P(5)(462),lamdaB => P(5)(494),lamdaOut => P(4)(462));
U_F5463: entity F port map(lamdaA => P(5)(463),lamdaB => P(5)(495),lamdaOut => P(4)(463));
U_F5464: entity F port map(lamdaA => P(5)(464),lamdaB => P(5)(496),lamdaOut => P(4)(464));
U_F5465: entity F port map(lamdaA => P(5)(465),lamdaB => P(5)(497),lamdaOut => P(4)(465));
U_F5466: entity F port map(lamdaA => P(5)(466),lamdaB => P(5)(498),lamdaOut => P(4)(466));
U_F5467: entity F port map(lamdaA => P(5)(467),lamdaB => P(5)(499),lamdaOut => P(4)(467));
U_F5468: entity F port map(lamdaA => P(5)(468),lamdaB => P(5)(500),lamdaOut => P(4)(468));
U_F5469: entity F port map(lamdaA => P(5)(469),lamdaB => P(5)(501),lamdaOut => P(4)(469));
U_F5470: entity F port map(lamdaA => P(5)(470),lamdaB => P(5)(502),lamdaOut => P(4)(470));
U_F5471: entity F port map(lamdaA => P(5)(471),lamdaB => P(5)(503),lamdaOut => P(4)(471));
U_F5472: entity F port map(lamdaA => P(5)(472),lamdaB => P(5)(504),lamdaOut => P(4)(472));
U_F5473: entity F port map(lamdaA => P(5)(473),lamdaB => P(5)(505),lamdaOut => P(4)(473));
U_F5474: entity F port map(lamdaA => P(5)(474),lamdaB => P(5)(506),lamdaOut => P(4)(474));
U_F5475: entity F port map(lamdaA => P(5)(475),lamdaB => P(5)(507),lamdaOut => P(4)(475));
U_F5476: entity F port map(lamdaA => P(5)(476),lamdaB => P(5)(508),lamdaOut => P(4)(476));
U_F5477: entity F port map(lamdaA => P(5)(477),lamdaB => P(5)(509),lamdaOut => P(4)(477));
U_F5478: entity F port map(lamdaA => P(5)(478),lamdaB => P(5)(510),lamdaOut => P(4)(478));
U_F5479: entity F port map(lamdaA => P(5)(479),lamdaB => P(5)(511),lamdaOut => P(4)(479));
U_G5480: entity G port map(lamdaA => P(5)(448),lamdaB => P(5)(480),s => s(5)(224),lamdaOut => P(4)(480));
U_G5481: entity G port map(lamdaA => P(5)(449),lamdaB => P(5)(481),s => s(5)(225),lamdaOut => P(4)(481));
U_G5482: entity G port map(lamdaA => P(5)(450),lamdaB => P(5)(482),s => s(5)(226),lamdaOut => P(4)(482));
U_G5483: entity G port map(lamdaA => P(5)(451),lamdaB => P(5)(483),s => s(5)(227),lamdaOut => P(4)(483));
U_G5484: entity G port map(lamdaA => P(5)(452),lamdaB => P(5)(484),s => s(5)(228),lamdaOut => P(4)(484));
U_G5485: entity G port map(lamdaA => P(5)(453),lamdaB => P(5)(485),s => s(5)(229),lamdaOut => P(4)(485));
U_G5486: entity G port map(lamdaA => P(5)(454),lamdaB => P(5)(486),s => s(5)(230),lamdaOut => P(4)(486));
U_G5487: entity G port map(lamdaA => P(5)(455),lamdaB => P(5)(487),s => s(5)(231),lamdaOut => P(4)(487));
U_G5488: entity G port map(lamdaA => P(5)(456),lamdaB => P(5)(488),s => s(5)(232),lamdaOut => P(4)(488));
U_G5489: entity G port map(lamdaA => P(5)(457),lamdaB => P(5)(489),s => s(5)(233),lamdaOut => P(4)(489));
U_G5490: entity G port map(lamdaA => P(5)(458),lamdaB => P(5)(490),s => s(5)(234),lamdaOut => P(4)(490));
U_G5491: entity G port map(lamdaA => P(5)(459),lamdaB => P(5)(491),s => s(5)(235),lamdaOut => P(4)(491));
U_G5492: entity G port map(lamdaA => P(5)(460),lamdaB => P(5)(492),s => s(5)(236),lamdaOut => P(4)(492));
U_G5493: entity G port map(lamdaA => P(5)(461),lamdaB => P(5)(493),s => s(5)(237),lamdaOut => P(4)(493));
U_G5494: entity G port map(lamdaA => P(5)(462),lamdaB => P(5)(494),s => s(5)(238),lamdaOut => P(4)(494));
U_G5495: entity G port map(lamdaA => P(5)(463),lamdaB => P(5)(495),s => s(5)(239),lamdaOut => P(4)(495));
U_G5496: entity G port map(lamdaA => P(5)(464),lamdaB => P(5)(496),s => s(5)(240),lamdaOut => P(4)(496));
U_G5497: entity G port map(lamdaA => P(5)(465),lamdaB => P(5)(497),s => s(5)(241),lamdaOut => P(4)(497));
U_G5498: entity G port map(lamdaA => P(5)(466),lamdaB => P(5)(498),s => s(5)(242),lamdaOut => P(4)(498));
U_G5499: entity G port map(lamdaA => P(5)(467),lamdaB => P(5)(499),s => s(5)(243),lamdaOut => P(4)(499));
U_G5500: entity G port map(lamdaA => P(5)(468),lamdaB => P(5)(500),s => s(5)(244),lamdaOut => P(4)(500));
U_G5501: entity G port map(lamdaA => P(5)(469),lamdaB => P(5)(501),s => s(5)(245),lamdaOut => P(4)(501));
U_G5502: entity G port map(lamdaA => P(5)(470),lamdaB => P(5)(502),s => s(5)(246),lamdaOut => P(4)(502));
U_G5503: entity G port map(lamdaA => P(5)(471),lamdaB => P(5)(503),s => s(5)(247),lamdaOut => P(4)(503));
U_G5504: entity G port map(lamdaA => P(5)(472),lamdaB => P(5)(504),s => s(5)(248),lamdaOut => P(4)(504));
U_G5505: entity G port map(lamdaA => P(5)(473),lamdaB => P(5)(505),s => s(5)(249),lamdaOut => P(4)(505));
U_G5506: entity G port map(lamdaA => P(5)(474),lamdaB => P(5)(506),s => s(5)(250),lamdaOut => P(4)(506));
U_G5507: entity G port map(lamdaA => P(5)(475),lamdaB => P(5)(507),s => s(5)(251),lamdaOut => P(4)(507));
U_G5508: entity G port map(lamdaA => P(5)(476),lamdaB => P(5)(508),s => s(5)(252),lamdaOut => P(4)(508));
U_G5509: entity G port map(lamdaA => P(5)(477),lamdaB => P(5)(509),s => s(5)(253),lamdaOut => P(4)(509));
U_G5510: entity G port map(lamdaA => P(5)(478),lamdaB => P(5)(510),s => s(5)(254),lamdaOut => P(4)(510));
U_G5511: entity G port map(lamdaA => P(5)(479),lamdaB => P(5)(511),s => s(5)(255),lamdaOut => P(4)(511));
U_F5512: entity F port map(lamdaA => P(5)(512),lamdaB => P(5)(544),lamdaOut => P(4)(512));
U_F5513: entity F port map(lamdaA => P(5)(513),lamdaB => P(5)(545),lamdaOut => P(4)(513));
U_F5514: entity F port map(lamdaA => P(5)(514),lamdaB => P(5)(546),lamdaOut => P(4)(514));
U_F5515: entity F port map(lamdaA => P(5)(515),lamdaB => P(5)(547),lamdaOut => P(4)(515));
U_F5516: entity F port map(lamdaA => P(5)(516),lamdaB => P(5)(548),lamdaOut => P(4)(516));
U_F5517: entity F port map(lamdaA => P(5)(517),lamdaB => P(5)(549),lamdaOut => P(4)(517));
U_F5518: entity F port map(lamdaA => P(5)(518),lamdaB => P(5)(550),lamdaOut => P(4)(518));
U_F5519: entity F port map(lamdaA => P(5)(519),lamdaB => P(5)(551),lamdaOut => P(4)(519));
U_F5520: entity F port map(lamdaA => P(5)(520),lamdaB => P(5)(552),lamdaOut => P(4)(520));
U_F5521: entity F port map(lamdaA => P(5)(521),lamdaB => P(5)(553),lamdaOut => P(4)(521));
U_F5522: entity F port map(lamdaA => P(5)(522),lamdaB => P(5)(554),lamdaOut => P(4)(522));
U_F5523: entity F port map(lamdaA => P(5)(523),lamdaB => P(5)(555),lamdaOut => P(4)(523));
U_F5524: entity F port map(lamdaA => P(5)(524),lamdaB => P(5)(556),lamdaOut => P(4)(524));
U_F5525: entity F port map(lamdaA => P(5)(525),lamdaB => P(5)(557),lamdaOut => P(4)(525));
U_F5526: entity F port map(lamdaA => P(5)(526),lamdaB => P(5)(558),lamdaOut => P(4)(526));
U_F5527: entity F port map(lamdaA => P(5)(527),lamdaB => P(5)(559),lamdaOut => P(4)(527));
U_F5528: entity F port map(lamdaA => P(5)(528),lamdaB => P(5)(560),lamdaOut => P(4)(528));
U_F5529: entity F port map(lamdaA => P(5)(529),lamdaB => P(5)(561),lamdaOut => P(4)(529));
U_F5530: entity F port map(lamdaA => P(5)(530),lamdaB => P(5)(562),lamdaOut => P(4)(530));
U_F5531: entity F port map(lamdaA => P(5)(531),lamdaB => P(5)(563),lamdaOut => P(4)(531));
U_F5532: entity F port map(lamdaA => P(5)(532),lamdaB => P(5)(564),lamdaOut => P(4)(532));
U_F5533: entity F port map(lamdaA => P(5)(533),lamdaB => P(5)(565),lamdaOut => P(4)(533));
U_F5534: entity F port map(lamdaA => P(5)(534),lamdaB => P(5)(566),lamdaOut => P(4)(534));
U_F5535: entity F port map(lamdaA => P(5)(535),lamdaB => P(5)(567),lamdaOut => P(4)(535));
U_F5536: entity F port map(lamdaA => P(5)(536),lamdaB => P(5)(568),lamdaOut => P(4)(536));
U_F5537: entity F port map(lamdaA => P(5)(537),lamdaB => P(5)(569),lamdaOut => P(4)(537));
U_F5538: entity F port map(lamdaA => P(5)(538),lamdaB => P(5)(570),lamdaOut => P(4)(538));
U_F5539: entity F port map(lamdaA => P(5)(539),lamdaB => P(5)(571),lamdaOut => P(4)(539));
U_F5540: entity F port map(lamdaA => P(5)(540),lamdaB => P(5)(572),lamdaOut => P(4)(540));
U_F5541: entity F port map(lamdaA => P(5)(541),lamdaB => P(5)(573),lamdaOut => P(4)(541));
U_F5542: entity F port map(lamdaA => P(5)(542),lamdaB => P(5)(574),lamdaOut => P(4)(542));
U_F5543: entity F port map(lamdaA => P(5)(543),lamdaB => P(5)(575),lamdaOut => P(4)(543));
U_G5544: entity G port map(lamdaA => P(5)(512),lamdaB => P(5)(544),s => s(5)(256),lamdaOut => P(4)(544));
U_G5545: entity G port map(lamdaA => P(5)(513),lamdaB => P(5)(545),s => s(5)(257),lamdaOut => P(4)(545));
U_G5546: entity G port map(lamdaA => P(5)(514),lamdaB => P(5)(546),s => s(5)(258),lamdaOut => P(4)(546));
U_G5547: entity G port map(lamdaA => P(5)(515),lamdaB => P(5)(547),s => s(5)(259),lamdaOut => P(4)(547));
U_G5548: entity G port map(lamdaA => P(5)(516),lamdaB => P(5)(548),s => s(5)(260),lamdaOut => P(4)(548));
U_G5549: entity G port map(lamdaA => P(5)(517),lamdaB => P(5)(549),s => s(5)(261),lamdaOut => P(4)(549));
U_G5550: entity G port map(lamdaA => P(5)(518),lamdaB => P(5)(550),s => s(5)(262),lamdaOut => P(4)(550));
U_G5551: entity G port map(lamdaA => P(5)(519),lamdaB => P(5)(551),s => s(5)(263),lamdaOut => P(4)(551));
U_G5552: entity G port map(lamdaA => P(5)(520),lamdaB => P(5)(552),s => s(5)(264),lamdaOut => P(4)(552));
U_G5553: entity G port map(lamdaA => P(5)(521),lamdaB => P(5)(553),s => s(5)(265),lamdaOut => P(4)(553));
U_G5554: entity G port map(lamdaA => P(5)(522),lamdaB => P(5)(554),s => s(5)(266),lamdaOut => P(4)(554));
U_G5555: entity G port map(lamdaA => P(5)(523),lamdaB => P(5)(555),s => s(5)(267),lamdaOut => P(4)(555));
U_G5556: entity G port map(lamdaA => P(5)(524),lamdaB => P(5)(556),s => s(5)(268),lamdaOut => P(4)(556));
U_G5557: entity G port map(lamdaA => P(5)(525),lamdaB => P(5)(557),s => s(5)(269),lamdaOut => P(4)(557));
U_G5558: entity G port map(lamdaA => P(5)(526),lamdaB => P(5)(558),s => s(5)(270),lamdaOut => P(4)(558));
U_G5559: entity G port map(lamdaA => P(5)(527),lamdaB => P(5)(559),s => s(5)(271),lamdaOut => P(4)(559));
U_G5560: entity G port map(lamdaA => P(5)(528),lamdaB => P(5)(560),s => s(5)(272),lamdaOut => P(4)(560));
U_G5561: entity G port map(lamdaA => P(5)(529),lamdaB => P(5)(561),s => s(5)(273),lamdaOut => P(4)(561));
U_G5562: entity G port map(lamdaA => P(5)(530),lamdaB => P(5)(562),s => s(5)(274),lamdaOut => P(4)(562));
U_G5563: entity G port map(lamdaA => P(5)(531),lamdaB => P(5)(563),s => s(5)(275),lamdaOut => P(4)(563));
U_G5564: entity G port map(lamdaA => P(5)(532),lamdaB => P(5)(564),s => s(5)(276),lamdaOut => P(4)(564));
U_G5565: entity G port map(lamdaA => P(5)(533),lamdaB => P(5)(565),s => s(5)(277),lamdaOut => P(4)(565));
U_G5566: entity G port map(lamdaA => P(5)(534),lamdaB => P(5)(566),s => s(5)(278),lamdaOut => P(4)(566));
U_G5567: entity G port map(lamdaA => P(5)(535),lamdaB => P(5)(567),s => s(5)(279),lamdaOut => P(4)(567));
U_G5568: entity G port map(lamdaA => P(5)(536),lamdaB => P(5)(568),s => s(5)(280),lamdaOut => P(4)(568));
U_G5569: entity G port map(lamdaA => P(5)(537),lamdaB => P(5)(569),s => s(5)(281),lamdaOut => P(4)(569));
U_G5570: entity G port map(lamdaA => P(5)(538),lamdaB => P(5)(570),s => s(5)(282),lamdaOut => P(4)(570));
U_G5571: entity G port map(lamdaA => P(5)(539),lamdaB => P(5)(571),s => s(5)(283),lamdaOut => P(4)(571));
U_G5572: entity G port map(lamdaA => P(5)(540),lamdaB => P(5)(572),s => s(5)(284),lamdaOut => P(4)(572));
U_G5573: entity G port map(lamdaA => P(5)(541),lamdaB => P(5)(573),s => s(5)(285),lamdaOut => P(4)(573));
U_G5574: entity G port map(lamdaA => P(5)(542),lamdaB => P(5)(574),s => s(5)(286),lamdaOut => P(4)(574));
U_G5575: entity G port map(lamdaA => P(5)(543),lamdaB => P(5)(575),s => s(5)(287),lamdaOut => P(4)(575));
U_F5576: entity F port map(lamdaA => P(5)(576),lamdaB => P(5)(608),lamdaOut => P(4)(576));
U_F5577: entity F port map(lamdaA => P(5)(577),lamdaB => P(5)(609),lamdaOut => P(4)(577));
U_F5578: entity F port map(lamdaA => P(5)(578),lamdaB => P(5)(610),lamdaOut => P(4)(578));
U_F5579: entity F port map(lamdaA => P(5)(579),lamdaB => P(5)(611),lamdaOut => P(4)(579));
U_F5580: entity F port map(lamdaA => P(5)(580),lamdaB => P(5)(612),lamdaOut => P(4)(580));
U_F5581: entity F port map(lamdaA => P(5)(581),lamdaB => P(5)(613),lamdaOut => P(4)(581));
U_F5582: entity F port map(lamdaA => P(5)(582),lamdaB => P(5)(614),lamdaOut => P(4)(582));
U_F5583: entity F port map(lamdaA => P(5)(583),lamdaB => P(5)(615),lamdaOut => P(4)(583));
U_F5584: entity F port map(lamdaA => P(5)(584),lamdaB => P(5)(616),lamdaOut => P(4)(584));
U_F5585: entity F port map(lamdaA => P(5)(585),lamdaB => P(5)(617),lamdaOut => P(4)(585));
U_F5586: entity F port map(lamdaA => P(5)(586),lamdaB => P(5)(618),lamdaOut => P(4)(586));
U_F5587: entity F port map(lamdaA => P(5)(587),lamdaB => P(5)(619),lamdaOut => P(4)(587));
U_F5588: entity F port map(lamdaA => P(5)(588),lamdaB => P(5)(620),lamdaOut => P(4)(588));
U_F5589: entity F port map(lamdaA => P(5)(589),lamdaB => P(5)(621),lamdaOut => P(4)(589));
U_F5590: entity F port map(lamdaA => P(5)(590),lamdaB => P(5)(622),lamdaOut => P(4)(590));
U_F5591: entity F port map(lamdaA => P(5)(591),lamdaB => P(5)(623),lamdaOut => P(4)(591));
U_F5592: entity F port map(lamdaA => P(5)(592),lamdaB => P(5)(624),lamdaOut => P(4)(592));
U_F5593: entity F port map(lamdaA => P(5)(593),lamdaB => P(5)(625),lamdaOut => P(4)(593));
U_F5594: entity F port map(lamdaA => P(5)(594),lamdaB => P(5)(626),lamdaOut => P(4)(594));
U_F5595: entity F port map(lamdaA => P(5)(595),lamdaB => P(5)(627),lamdaOut => P(4)(595));
U_F5596: entity F port map(lamdaA => P(5)(596),lamdaB => P(5)(628),lamdaOut => P(4)(596));
U_F5597: entity F port map(lamdaA => P(5)(597),lamdaB => P(5)(629),lamdaOut => P(4)(597));
U_F5598: entity F port map(lamdaA => P(5)(598),lamdaB => P(5)(630),lamdaOut => P(4)(598));
U_F5599: entity F port map(lamdaA => P(5)(599),lamdaB => P(5)(631),lamdaOut => P(4)(599));
U_F5600: entity F port map(lamdaA => P(5)(600),lamdaB => P(5)(632),lamdaOut => P(4)(600));
U_F5601: entity F port map(lamdaA => P(5)(601),lamdaB => P(5)(633),lamdaOut => P(4)(601));
U_F5602: entity F port map(lamdaA => P(5)(602),lamdaB => P(5)(634),lamdaOut => P(4)(602));
U_F5603: entity F port map(lamdaA => P(5)(603),lamdaB => P(5)(635),lamdaOut => P(4)(603));
U_F5604: entity F port map(lamdaA => P(5)(604),lamdaB => P(5)(636),lamdaOut => P(4)(604));
U_F5605: entity F port map(lamdaA => P(5)(605),lamdaB => P(5)(637),lamdaOut => P(4)(605));
U_F5606: entity F port map(lamdaA => P(5)(606),lamdaB => P(5)(638),lamdaOut => P(4)(606));
U_F5607: entity F port map(lamdaA => P(5)(607),lamdaB => P(5)(639),lamdaOut => P(4)(607));
U_G5608: entity G port map(lamdaA => P(5)(576),lamdaB => P(5)(608),s => s(5)(288),lamdaOut => P(4)(608));
U_G5609: entity G port map(lamdaA => P(5)(577),lamdaB => P(5)(609),s => s(5)(289),lamdaOut => P(4)(609));
U_G5610: entity G port map(lamdaA => P(5)(578),lamdaB => P(5)(610),s => s(5)(290),lamdaOut => P(4)(610));
U_G5611: entity G port map(lamdaA => P(5)(579),lamdaB => P(5)(611),s => s(5)(291),lamdaOut => P(4)(611));
U_G5612: entity G port map(lamdaA => P(5)(580),lamdaB => P(5)(612),s => s(5)(292),lamdaOut => P(4)(612));
U_G5613: entity G port map(lamdaA => P(5)(581),lamdaB => P(5)(613),s => s(5)(293),lamdaOut => P(4)(613));
U_G5614: entity G port map(lamdaA => P(5)(582),lamdaB => P(5)(614),s => s(5)(294),lamdaOut => P(4)(614));
U_G5615: entity G port map(lamdaA => P(5)(583),lamdaB => P(5)(615),s => s(5)(295),lamdaOut => P(4)(615));
U_G5616: entity G port map(lamdaA => P(5)(584),lamdaB => P(5)(616),s => s(5)(296),lamdaOut => P(4)(616));
U_G5617: entity G port map(lamdaA => P(5)(585),lamdaB => P(5)(617),s => s(5)(297),lamdaOut => P(4)(617));
U_G5618: entity G port map(lamdaA => P(5)(586),lamdaB => P(5)(618),s => s(5)(298),lamdaOut => P(4)(618));
U_G5619: entity G port map(lamdaA => P(5)(587),lamdaB => P(5)(619),s => s(5)(299),lamdaOut => P(4)(619));
U_G5620: entity G port map(lamdaA => P(5)(588),lamdaB => P(5)(620),s => s(5)(300),lamdaOut => P(4)(620));
U_G5621: entity G port map(lamdaA => P(5)(589),lamdaB => P(5)(621),s => s(5)(301),lamdaOut => P(4)(621));
U_G5622: entity G port map(lamdaA => P(5)(590),lamdaB => P(5)(622),s => s(5)(302),lamdaOut => P(4)(622));
U_G5623: entity G port map(lamdaA => P(5)(591),lamdaB => P(5)(623),s => s(5)(303),lamdaOut => P(4)(623));
U_G5624: entity G port map(lamdaA => P(5)(592),lamdaB => P(5)(624),s => s(5)(304),lamdaOut => P(4)(624));
U_G5625: entity G port map(lamdaA => P(5)(593),lamdaB => P(5)(625),s => s(5)(305),lamdaOut => P(4)(625));
U_G5626: entity G port map(lamdaA => P(5)(594),lamdaB => P(5)(626),s => s(5)(306),lamdaOut => P(4)(626));
U_G5627: entity G port map(lamdaA => P(5)(595),lamdaB => P(5)(627),s => s(5)(307),lamdaOut => P(4)(627));
U_G5628: entity G port map(lamdaA => P(5)(596),lamdaB => P(5)(628),s => s(5)(308),lamdaOut => P(4)(628));
U_G5629: entity G port map(lamdaA => P(5)(597),lamdaB => P(5)(629),s => s(5)(309),lamdaOut => P(4)(629));
U_G5630: entity G port map(lamdaA => P(5)(598),lamdaB => P(5)(630),s => s(5)(310),lamdaOut => P(4)(630));
U_G5631: entity G port map(lamdaA => P(5)(599),lamdaB => P(5)(631),s => s(5)(311),lamdaOut => P(4)(631));
U_G5632: entity G port map(lamdaA => P(5)(600),lamdaB => P(5)(632),s => s(5)(312),lamdaOut => P(4)(632));
U_G5633: entity G port map(lamdaA => P(5)(601),lamdaB => P(5)(633),s => s(5)(313),lamdaOut => P(4)(633));
U_G5634: entity G port map(lamdaA => P(5)(602),lamdaB => P(5)(634),s => s(5)(314),lamdaOut => P(4)(634));
U_G5635: entity G port map(lamdaA => P(5)(603),lamdaB => P(5)(635),s => s(5)(315),lamdaOut => P(4)(635));
U_G5636: entity G port map(lamdaA => P(5)(604),lamdaB => P(5)(636),s => s(5)(316),lamdaOut => P(4)(636));
U_G5637: entity G port map(lamdaA => P(5)(605),lamdaB => P(5)(637),s => s(5)(317),lamdaOut => P(4)(637));
U_G5638: entity G port map(lamdaA => P(5)(606),lamdaB => P(5)(638),s => s(5)(318),lamdaOut => P(4)(638));
U_G5639: entity G port map(lamdaA => P(5)(607),lamdaB => P(5)(639),s => s(5)(319),lamdaOut => P(4)(639));
U_F5640: entity F port map(lamdaA => P(5)(640),lamdaB => P(5)(672),lamdaOut => P(4)(640));
U_F5641: entity F port map(lamdaA => P(5)(641),lamdaB => P(5)(673),lamdaOut => P(4)(641));
U_F5642: entity F port map(lamdaA => P(5)(642),lamdaB => P(5)(674),lamdaOut => P(4)(642));
U_F5643: entity F port map(lamdaA => P(5)(643),lamdaB => P(5)(675),lamdaOut => P(4)(643));
U_F5644: entity F port map(lamdaA => P(5)(644),lamdaB => P(5)(676),lamdaOut => P(4)(644));
U_F5645: entity F port map(lamdaA => P(5)(645),lamdaB => P(5)(677),lamdaOut => P(4)(645));
U_F5646: entity F port map(lamdaA => P(5)(646),lamdaB => P(5)(678),lamdaOut => P(4)(646));
U_F5647: entity F port map(lamdaA => P(5)(647),lamdaB => P(5)(679),lamdaOut => P(4)(647));
U_F5648: entity F port map(lamdaA => P(5)(648),lamdaB => P(5)(680),lamdaOut => P(4)(648));
U_F5649: entity F port map(lamdaA => P(5)(649),lamdaB => P(5)(681),lamdaOut => P(4)(649));
U_F5650: entity F port map(lamdaA => P(5)(650),lamdaB => P(5)(682),lamdaOut => P(4)(650));
U_F5651: entity F port map(lamdaA => P(5)(651),lamdaB => P(5)(683),lamdaOut => P(4)(651));
U_F5652: entity F port map(lamdaA => P(5)(652),lamdaB => P(5)(684),lamdaOut => P(4)(652));
U_F5653: entity F port map(lamdaA => P(5)(653),lamdaB => P(5)(685),lamdaOut => P(4)(653));
U_F5654: entity F port map(lamdaA => P(5)(654),lamdaB => P(5)(686),lamdaOut => P(4)(654));
U_F5655: entity F port map(lamdaA => P(5)(655),lamdaB => P(5)(687),lamdaOut => P(4)(655));
U_F5656: entity F port map(lamdaA => P(5)(656),lamdaB => P(5)(688),lamdaOut => P(4)(656));
U_F5657: entity F port map(lamdaA => P(5)(657),lamdaB => P(5)(689),lamdaOut => P(4)(657));
U_F5658: entity F port map(lamdaA => P(5)(658),lamdaB => P(5)(690),lamdaOut => P(4)(658));
U_F5659: entity F port map(lamdaA => P(5)(659),lamdaB => P(5)(691),lamdaOut => P(4)(659));
U_F5660: entity F port map(lamdaA => P(5)(660),lamdaB => P(5)(692),lamdaOut => P(4)(660));
U_F5661: entity F port map(lamdaA => P(5)(661),lamdaB => P(5)(693),lamdaOut => P(4)(661));
U_F5662: entity F port map(lamdaA => P(5)(662),lamdaB => P(5)(694),lamdaOut => P(4)(662));
U_F5663: entity F port map(lamdaA => P(5)(663),lamdaB => P(5)(695),lamdaOut => P(4)(663));
U_F5664: entity F port map(lamdaA => P(5)(664),lamdaB => P(5)(696),lamdaOut => P(4)(664));
U_F5665: entity F port map(lamdaA => P(5)(665),lamdaB => P(5)(697),lamdaOut => P(4)(665));
U_F5666: entity F port map(lamdaA => P(5)(666),lamdaB => P(5)(698),lamdaOut => P(4)(666));
U_F5667: entity F port map(lamdaA => P(5)(667),lamdaB => P(5)(699),lamdaOut => P(4)(667));
U_F5668: entity F port map(lamdaA => P(5)(668),lamdaB => P(5)(700),lamdaOut => P(4)(668));
U_F5669: entity F port map(lamdaA => P(5)(669),lamdaB => P(5)(701),lamdaOut => P(4)(669));
U_F5670: entity F port map(lamdaA => P(5)(670),lamdaB => P(5)(702),lamdaOut => P(4)(670));
U_F5671: entity F port map(lamdaA => P(5)(671),lamdaB => P(5)(703),lamdaOut => P(4)(671));
U_G5672: entity G port map(lamdaA => P(5)(640),lamdaB => P(5)(672),s => s(5)(320),lamdaOut => P(4)(672));
U_G5673: entity G port map(lamdaA => P(5)(641),lamdaB => P(5)(673),s => s(5)(321),lamdaOut => P(4)(673));
U_G5674: entity G port map(lamdaA => P(5)(642),lamdaB => P(5)(674),s => s(5)(322),lamdaOut => P(4)(674));
U_G5675: entity G port map(lamdaA => P(5)(643),lamdaB => P(5)(675),s => s(5)(323),lamdaOut => P(4)(675));
U_G5676: entity G port map(lamdaA => P(5)(644),lamdaB => P(5)(676),s => s(5)(324),lamdaOut => P(4)(676));
U_G5677: entity G port map(lamdaA => P(5)(645),lamdaB => P(5)(677),s => s(5)(325),lamdaOut => P(4)(677));
U_G5678: entity G port map(lamdaA => P(5)(646),lamdaB => P(5)(678),s => s(5)(326),lamdaOut => P(4)(678));
U_G5679: entity G port map(lamdaA => P(5)(647),lamdaB => P(5)(679),s => s(5)(327),lamdaOut => P(4)(679));
U_G5680: entity G port map(lamdaA => P(5)(648),lamdaB => P(5)(680),s => s(5)(328),lamdaOut => P(4)(680));
U_G5681: entity G port map(lamdaA => P(5)(649),lamdaB => P(5)(681),s => s(5)(329),lamdaOut => P(4)(681));
U_G5682: entity G port map(lamdaA => P(5)(650),lamdaB => P(5)(682),s => s(5)(330),lamdaOut => P(4)(682));
U_G5683: entity G port map(lamdaA => P(5)(651),lamdaB => P(5)(683),s => s(5)(331),lamdaOut => P(4)(683));
U_G5684: entity G port map(lamdaA => P(5)(652),lamdaB => P(5)(684),s => s(5)(332),lamdaOut => P(4)(684));
U_G5685: entity G port map(lamdaA => P(5)(653),lamdaB => P(5)(685),s => s(5)(333),lamdaOut => P(4)(685));
U_G5686: entity G port map(lamdaA => P(5)(654),lamdaB => P(5)(686),s => s(5)(334),lamdaOut => P(4)(686));
U_G5687: entity G port map(lamdaA => P(5)(655),lamdaB => P(5)(687),s => s(5)(335),lamdaOut => P(4)(687));
U_G5688: entity G port map(lamdaA => P(5)(656),lamdaB => P(5)(688),s => s(5)(336),lamdaOut => P(4)(688));
U_G5689: entity G port map(lamdaA => P(5)(657),lamdaB => P(5)(689),s => s(5)(337),lamdaOut => P(4)(689));
U_G5690: entity G port map(lamdaA => P(5)(658),lamdaB => P(5)(690),s => s(5)(338),lamdaOut => P(4)(690));
U_G5691: entity G port map(lamdaA => P(5)(659),lamdaB => P(5)(691),s => s(5)(339),lamdaOut => P(4)(691));
U_G5692: entity G port map(lamdaA => P(5)(660),lamdaB => P(5)(692),s => s(5)(340),lamdaOut => P(4)(692));
U_G5693: entity G port map(lamdaA => P(5)(661),lamdaB => P(5)(693),s => s(5)(341),lamdaOut => P(4)(693));
U_G5694: entity G port map(lamdaA => P(5)(662),lamdaB => P(5)(694),s => s(5)(342),lamdaOut => P(4)(694));
U_G5695: entity G port map(lamdaA => P(5)(663),lamdaB => P(5)(695),s => s(5)(343),lamdaOut => P(4)(695));
U_G5696: entity G port map(lamdaA => P(5)(664),lamdaB => P(5)(696),s => s(5)(344),lamdaOut => P(4)(696));
U_G5697: entity G port map(lamdaA => P(5)(665),lamdaB => P(5)(697),s => s(5)(345),lamdaOut => P(4)(697));
U_G5698: entity G port map(lamdaA => P(5)(666),lamdaB => P(5)(698),s => s(5)(346),lamdaOut => P(4)(698));
U_G5699: entity G port map(lamdaA => P(5)(667),lamdaB => P(5)(699),s => s(5)(347),lamdaOut => P(4)(699));
U_G5700: entity G port map(lamdaA => P(5)(668),lamdaB => P(5)(700),s => s(5)(348),lamdaOut => P(4)(700));
U_G5701: entity G port map(lamdaA => P(5)(669),lamdaB => P(5)(701),s => s(5)(349),lamdaOut => P(4)(701));
U_G5702: entity G port map(lamdaA => P(5)(670),lamdaB => P(5)(702),s => s(5)(350),lamdaOut => P(4)(702));
U_G5703: entity G port map(lamdaA => P(5)(671),lamdaB => P(5)(703),s => s(5)(351),lamdaOut => P(4)(703));
U_F5704: entity F port map(lamdaA => P(5)(704),lamdaB => P(5)(736),lamdaOut => P(4)(704));
U_F5705: entity F port map(lamdaA => P(5)(705),lamdaB => P(5)(737),lamdaOut => P(4)(705));
U_F5706: entity F port map(lamdaA => P(5)(706),lamdaB => P(5)(738),lamdaOut => P(4)(706));
U_F5707: entity F port map(lamdaA => P(5)(707),lamdaB => P(5)(739),lamdaOut => P(4)(707));
U_F5708: entity F port map(lamdaA => P(5)(708),lamdaB => P(5)(740),lamdaOut => P(4)(708));
U_F5709: entity F port map(lamdaA => P(5)(709),lamdaB => P(5)(741),lamdaOut => P(4)(709));
U_F5710: entity F port map(lamdaA => P(5)(710),lamdaB => P(5)(742),lamdaOut => P(4)(710));
U_F5711: entity F port map(lamdaA => P(5)(711),lamdaB => P(5)(743),lamdaOut => P(4)(711));
U_F5712: entity F port map(lamdaA => P(5)(712),lamdaB => P(5)(744),lamdaOut => P(4)(712));
U_F5713: entity F port map(lamdaA => P(5)(713),lamdaB => P(5)(745),lamdaOut => P(4)(713));
U_F5714: entity F port map(lamdaA => P(5)(714),lamdaB => P(5)(746),lamdaOut => P(4)(714));
U_F5715: entity F port map(lamdaA => P(5)(715),lamdaB => P(5)(747),lamdaOut => P(4)(715));
U_F5716: entity F port map(lamdaA => P(5)(716),lamdaB => P(5)(748),lamdaOut => P(4)(716));
U_F5717: entity F port map(lamdaA => P(5)(717),lamdaB => P(5)(749),lamdaOut => P(4)(717));
U_F5718: entity F port map(lamdaA => P(5)(718),lamdaB => P(5)(750),lamdaOut => P(4)(718));
U_F5719: entity F port map(lamdaA => P(5)(719),lamdaB => P(5)(751),lamdaOut => P(4)(719));
U_F5720: entity F port map(lamdaA => P(5)(720),lamdaB => P(5)(752),lamdaOut => P(4)(720));
U_F5721: entity F port map(lamdaA => P(5)(721),lamdaB => P(5)(753),lamdaOut => P(4)(721));
U_F5722: entity F port map(lamdaA => P(5)(722),lamdaB => P(5)(754),lamdaOut => P(4)(722));
U_F5723: entity F port map(lamdaA => P(5)(723),lamdaB => P(5)(755),lamdaOut => P(4)(723));
U_F5724: entity F port map(lamdaA => P(5)(724),lamdaB => P(5)(756),lamdaOut => P(4)(724));
U_F5725: entity F port map(lamdaA => P(5)(725),lamdaB => P(5)(757),lamdaOut => P(4)(725));
U_F5726: entity F port map(lamdaA => P(5)(726),lamdaB => P(5)(758),lamdaOut => P(4)(726));
U_F5727: entity F port map(lamdaA => P(5)(727),lamdaB => P(5)(759),lamdaOut => P(4)(727));
U_F5728: entity F port map(lamdaA => P(5)(728),lamdaB => P(5)(760),lamdaOut => P(4)(728));
U_F5729: entity F port map(lamdaA => P(5)(729),lamdaB => P(5)(761),lamdaOut => P(4)(729));
U_F5730: entity F port map(lamdaA => P(5)(730),lamdaB => P(5)(762),lamdaOut => P(4)(730));
U_F5731: entity F port map(lamdaA => P(5)(731),lamdaB => P(5)(763),lamdaOut => P(4)(731));
U_F5732: entity F port map(lamdaA => P(5)(732),lamdaB => P(5)(764),lamdaOut => P(4)(732));
U_F5733: entity F port map(lamdaA => P(5)(733),lamdaB => P(5)(765),lamdaOut => P(4)(733));
U_F5734: entity F port map(lamdaA => P(5)(734),lamdaB => P(5)(766),lamdaOut => P(4)(734));
U_F5735: entity F port map(lamdaA => P(5)(735),lamdaB => P(5)(767),lamdaOut => P(4)(735));
U_G5736: entity G port map(lamdaA => P(5)(704),lamdaB => P(5)(736),s => s(5)(352),lamdaOut => P(4)(736));
U_G5737: entity G port map(lamdaA => P(5)(705),lamdaB => P(5)(737),s => s(5)(353),lamdaOut => P(4)(737));
U_G5738: entity G port map(lamdaA => P(5)(706),lamdaB => P(5)(738),s => s(5)(354),lamdaOut => P(4)(738));
U_G5739: entity G port map(lamdaA => P(5)(707),lamdaB => P(5)(739),s => s(5)(355),lamdaOut => P(4)(739));
U_G5740: entity G port map(lamdaA => P(5)(708),lamdaB => P(5)(740),s => s(5)(356),lamdaOut => P(4)(740));
U_G5741: entity G port map(lamdaA => P(5)(709),lamdaB => P(5)(741),s => s(5)(357),lamdaOut => P(4)(741));
U_G5742: entity G port map(lamdaA => P(5)(710),lamdaB => P(5)(742),s => s(5)(358),lamdaOut => P(4)(742));
U_G5743: entity G port map(lamdaA => P(5)(711),lamdaB => P(5)(743),s => s(5)(359),lamdaOut => P(4)(743));
U_G5744: entity G port map(lamdaA => P(5)(712),lamdaB => P(5)(744),s => s(5)(360),lamdaOut => P(4)(744));
U_G5745: entity G port map(lamdaA => P(5)(713),lamdaB => P(5)(745),s => s(5)(361),lamdaOut => P(4)(745));
U_G5746: entity G port map(lamdaA => P(5)(714),lamdaB => P(5)(746),s => s(5)(362),lamdaOut => P(4)(746));
U_G5747: entity G port map(lamdaA => P(5)(715),lamdaB => P(5)(747),s => s(5)(363),lamdaOut => P(4)(747));
U_G5748: entity G port map(lamdaA => P(5)(716),lamdaB => P(5)(748),s => s(5)(364),lamdaOut => P(4)(748));
U_G5749: entity G port map(lamdaA => P(5)(717),lamdaB => P(5)(749),s => s(5)(365),lamdaOut => P(4)(749));
U_G5750: entity G port map(lamdaA => P(5)(718),lamdaB => P(5)(750),s => s(5)(366),lamdaOut => P(4)(750));
U_G5751: entity G port map(lamdaA => P(5)(719),lamdaB => P(5)(751),s => s(5)(367),lamdaOut => P(4)(751));
U_G5752: entity G port map(lamdaA => P(5)(720),lamdaB => P(5)(752),s => s(5)(368),lamdaOut => P(4)(752));
U_G5753: entity G port map(lamdaA => P(5)(721),lamdaB => P(5)(753),s => s(5)(369),lamdaOut => P(4)(753));
U_G5754: entity G port map(lamdaA => P(5)(722),lamdaB => P(5)(754),s => s(5)(370),lamdaOut => P(4)(754));
U_G5755: entity G port map(lamdaA => P(5)(723),lamdaB => P(5)(755),s => s(5)(371),lamdaOut => P(4)(755));
U_G5756: entity G port map(lamdaA => P(5)(724),lamdaB => P(5)(756),s => s(5)(372),lamdaOut => P(4)(756));
U_G5757: entity G port map(lamdaA => P(5)(725),lamdaB => P(5)(757),s => s(5)(373),lamdaOut => P(4)(757));
U_G5758: entity G port map(lamdaA => P(5)(726),lamdaB => P(5)(758),s => s(5)(374),lamdaOut => P(4)(758));
U_G5759: entity G port map(lamdaA => P(5)(727),lamdaB => P(5)(759),s => s(5)(375),lamdaOut => P(4)(759));
U_G5760: entity G port map(lamdaA => P(5)(728),lamdaB => P(5)(760),s => s(5)(376),lamdaOut => P(4)(760));
U_G5761: entity G port map(lamdaA => P(5)(729),lamdaB => P(5)(761),s => s(5)(377),lamdaOut => P(4)(761));
U_G5762: entity G port map(lamdaA => P(5)(730),lamdaB => P(5)(762),s => s(5)(378),lamdaOut => P(4)(762));
U_G5763: entity G port map(lamdaA => P(5)(731),lamdaB => P(5)(763),s => s(5)(379),lamdaOut => P(4)(763));
U_G5764: entity G port map(lamdaA => P(5)(732),lamdaB => P(5)(764),s => s(5)(380),lamdaOut => P(4)(764));
U_G5765: entity G port map(lamdaA => P(5)(733),lamdaB => P(5)(765),s => s(5)(381),lamdaOut => P(4)(765));
U_G5766: entity G port map(lamdaA => P(5)(734),lamdaB => P(5)(766),s => s(5)(382),lamdaOut => P(4)(766));
U_G5767: entity G port map(lamdaA => P(5)(735),lamdaB => P(5)(767),s => s(5)(383),lamdaOut => P(4)(767));
U_F5768: entity F port map(lamdaA => P(5)(768),lamdaB => P(5)(800),lamdaOut => P(4)(768));
U_F5769: entity F port map(lamdaA => P(5)(769),lamdaB => P(5)(801),lamdaOut => P(4)(769));
U_F5770: entity F port map(lamdaA => P(5)(770),lamdaB => P(5)(802),lamdaOut => P(4)(770));
U_F5771: entity F port map(lamdaA => P(5)(771),lamdaB => P(5)(803),lamdaOut => P(4)(771));
U_F5772: entity F port map(lamdaA => P(5)(772),lamdaB => P(5)(804),lamdaOut => P(4)(772));
U_F5773: entity F port map(lamdaA => P(5)(773),lamdaB => P(5)(805),lamdaOut => P(4)(773));
U_F5774: entity F port map(lamdaA => P(5)(774),lamdaB => P(5)(806),lamdaOut => P(4)(774));
U_F5775: entity F port map(lamdaA => P(5)(775),lamdaB => P(5)(807),lamdaOut => P(4)(775));
U_F5776: entity F port map(lamdaA => P(5)(776),lamdaB => P(5)(808),lamdaOut => P(4)(776));
U_F5777: entity F port map(lamdaA => P(5)(777),lamdaB => P(5)(809),lamdaOut => P(4)(777));
U_F5778: entity F port map(lamdaA => P(5)(778),lamdaB => P(5)(810),lamdaOut => P(4)(778));
U_F5779: entity F port map(lamdaA => P(5)(779),lamdaB => P(5)(811),lamdaOut => P(4)(779));
U_F5780: entity F port map(lamdaA => P(5)(780),lamdaB => P(5)(812),lamdaOut => P(4)(780));
U_F5781: entity F port map(lamdaA => P(5)(781),lamdaB => P(5)(813),lamdaOut => P(4)(781));
U_F5782: entity F port map(lamdaA => P(5)(782),lamdaB => P(5)(814),lamdaOut => P(4)(782));
U_F5783: entity F port map(lamdaA => P(5)(783),lamdaB => P(5)(815),lamdaOut => P(4)(783));
U_F5784: entity F port map(lamdaA => P(5)(784),lamdaB => P(5)(816),lamdaOut => P(4)(784));
U_F5785: entity F port map(lamdaA => P(5)(785),lamdaB => P(5)(817),lamdaOut => P(4)(785));
U_F5786: entity F port map(lamdaA => P(5)(786),lamdaB => P(5)(818),lamdaOut => P(4)(786));
U_F5787: entity F port map(lamdaA => P(5)(787),lamdaB => P(5)(819),lamdaOut => P(4)(787));
U_F5788: entity F port map(lamdaA => P(5)(788),lamdaB => P(5)(820),lamdaOut => P(4)(788));
U_F5789: entity F port map(lamdaA => P(5)(789),lamdaB => P(5)(821),lamdaOut => P(4)(789));
U_F5790: entity F port map(lamdaA => P(5)(790),lamdaB => P(5)(822),lamdaOut => P(4)(790));
U_F5791: entity F port map(lamdaA => P(5)(791),lamdaB => P(5)(823),lamdaOut => P(4)(791));
U_F5792: entity F port map(lamdaA => P(5)(792),lamdaB => P(5)(824),lamdaOut => P(4)(792));
U_F5793: entity F port map(lamdaA => P(5)(793),lamdaB => P(5)(825),lamdaOut => P(4)(793));
U_F5794: entity F port map(lamdaA => P(5)(794),lamdaB => P(5)(826),lamdaOut => P(4)(794));
U_F5795: entity F port map(lamdaA => P(5)(795),lamdaB => P(5)(827),lamdaOut => P(4)(795));
U_F5796: entity F port map(lamdaA => P(5)(796),lamdaB => P(5)(828),lamdaOut => P(4)(796));
U_F5797: entity F port map(lamdaA => P(5)(797),lamdaB => P(5)(829),lamdaOut => P(4)(797));
U_F5798: entity F port map(lamdaA => P(5)(798),lamdaB => P(5)(830),lamdaOut => P(4)(798));
U_F5799: entity F port map(lamdaA => P(5)(799),lamdaB => P(5)(831),lamdaOut => P(4)(799));
U_G5800: entity G port map(lamdaA => P(5)(768),lamdaB => P(5)(800),s => s(5)(384),lamdaOut => P(4)(800));
U_G5801: entity G port map(lamdaA => P(5)(769),lamdaB => P(5)(801),s => s(5)(385),lamdaOut => P(4)(801));
U_G5802: entity G port map(lamdaA => P(5)(770),lamdaB => P(5)(802),s => s(5)(386),lamdaOut => P(4)(802));
U_G5803: entity G port map(lamdaA => P(5)(771),lamdaB => P(5)(803),s => s(5)(387),lamdaOut => P(4)(803));
U_G5804: entity G port map(lamdaA => P(5)(772),lamdaB => P(5)(804),s => s(5)(388),lamdaOut => P(4)(804));
U_G5805: entity G port map(lamdaA => P(5)(773),lamdaB => P(5)(805),s => s(5)(389),lamdaOut => P(4)(805));
U_G5806: entity G port map(lamdaA => P(5)(774),lamdaB => P(5)(806),s => s(5)(390),lamdaOut => P(4)(806));
U_G5807: entity G port map(lamdaA => P(5)(775),lamdaB => P(5)(807),s => s(5)(391),lamdaOut => P(4)(807));
U_G5808: entity G port map(lamdaA => P(5)(776),lamdaB => P(5)(808),s => s(5)(392),lamdaOut => P(4)(808));
U_G5809: entity G port map(lamdaA => P(5)(777),lamdaB => P(5)(809),s => s(5)(393),lamdaOut => P(4)(809));
U_G5810: entity G port map(lamdaA => P(5)(778),lamdaB => P(5)(810),s => s(5)(394),lamdaOut => P(4)(810));
U_G5811: entity G port map(lamdaA => P(5)(779),lamdaB => P(5)(811),s => s(5)(395),lamdaOut => P(4)(811));
U_G5812: entity G port map(lamdaA => P(5)(780),lamdaB => P(5)(812),s => s(5)(396),lamdaOut => P(4)(812));
U_G5813: entity G port map(lamdaA => P(5)(781),lamdaB => P(5)(813),s => s(5)(397),lamdaOut => P(4)(813));
U_G5814: entity G port map(lamdaA => P(5)(782),lamdaB => P(5)(814),s => s(5)(398),lamdaOut => P(4)(814));
U_G5815: entity G port map(lamdaA => P(5)(783),lamdaB => P(5)(815),s => s(5)(399),lamdaOut => P(4)(815));
U_G5816: entity G port map(lamdaA => P(5)(784),lamdaB => P(5)(816),s => s(5)(400),lamdaOut => P(4)(816));
U_G5817: entity G port map(lamdaA => P(5)(785),lamdaB => P(5)(817),s => s(5)(401),lamdaOut => P(4)(817));
U_G5818: entity G port map(lamdaA => P(5)(786),lamdaB => P(5)(818),s => s(5)(402),lamdaOut => P(4)(818));
U_G5819: entity G port map(lamdaA => P(5)(787),lamdaB => P(5)(819),s => s(5)(403),lamdaOut => P(4)(819));
U_G5820: entity G port map(lamdaA => P(5)(788),lamdaB => P(5)(820),s => s(5)(404),lamdaOut => P(4)(820));
U_G5821: entity G port map(lamdaA => P(5)(789),lamdaB => P(5)(821),s => s(5)(405),lamdaOut => P(4)(821));
U_G5822: entity G port map(lamdaA => P(5)(790),lamdaB => P(5)(822),s => s(5)(406),lamdaOut => P(4)(822));
U_G5823: entity G port map(lamdaA => P(5)(791),lamdaB => P(5)(823),s => s(5)(407),lamdaOut => P(4)(823));
U_G5824: entity G port map(lamdaA => P(5)(792),lamdaB => P(5)(824),s => s(5)(408),lamdaOut => P(4)(824));
U_G5825: entity G port map(lamdaA => P(5)(793),lamdaB => P(5)(825),s => s(5)(409),lamdaOut => P(4)(825));
U_G5826: entity G port map(lamdaA => P(5)(794),lamdaB => P(5)(826),s => s(5)(410),lamdaOut => P(4)(826));
U_G5827: entity G port map(lamdaA => P(5)(795),lamdaB => P(5)(827),s => s(5)(411),lamdaOut => P(4)(827));
U_G5828: entity G port map(lamdaA => P(5)(796),lamdaB => P(5)(828),s => s(5)(412),lamdaOut => P(4)(828));
U_G5829: entity G port map(lamdaA => P(5)(797),lamdaB => P(5)(829),s => s(5)(413),lamdaOut => P(4)(829));
U_G5830: entity G port map(lamdaA => P(5)(798),lamdaB => P(5)(830),s => s(5)(414),lamdaOut => P(4)(830));
U_G5831: entity G port map(lamdaA => P(5)(799),lamdaB => P(5)(831),s => s(5)(415),lamdaOut => P(4)(831));
U_F5832: entity F port map(lamdaA => P(5)(832),lamdaB => P(5)(864),lamdaOut => P(4)(832));
U_F5833: entity F port map(lamdaA => P(5)(833),lamdaB => P(5)(865),lamdaOut => P(4)(833));
U_F5834: entity F port map(lamdaA => P(5)(834),lamdaB => P(5)(866),lamdaOut => P(4)(834));
U_F5835: entity F port map(lamdaA => P(5)(835),lamdaB => P(5)(867),lamdaOut => P(4)(835));
U_F5836: entity F port map(lamdaA => P(5)(836),lamdaB => P(5)(868),lamdaOut => P(4)(836));
U_F5837: entity F port map(lamdaA => P(5)(837),lamdaB => P(5)(869),lamdaOut => P(4)(837));
U_F5838: entity F port map(lamdaA => P(5)(838),lamdaB => P(5)(870),lamdaOut => P(4)(838));
U_F5839: entity F port map(lamdaA => P(5)(839),lamdaB => P(5)(871),lamdaOut => P(4)(839));
U_F5840: entity F port map(lamdaA => P(5)(840),lamdaB => P(5)(872),lamdaOut => P(4)(840));
U_F5841: entity F port map(lamdaA => P(5)(841),lamdaB => P(5)(873),lamdaOut => P(4)(841));
U_F5842: entity F port map(lamdaA => P(5)(842),lamdaB => P(5)(874),lamdaOut => P(4)(842));
U_F5843: entity F port map(lamdaA => P(5)(843),lamdaB => P(5)(875),lamdaOut => P(4)(843));
U_F5844: entity F port map(lamdaA => P(5)(844),lamdaB => P(5)(876),lamdaOut => P(4)(844));
U_F5845: entity F port map(lamdaA => P(5)(845),lamdaB => P(5)(877),lamdaOut => P(4)(845));
U_F5846: entity F port map(lamdaA => P(5)(846),lamdaB => P(5)(878),lamdaOut => P(4)(846));
U_F5847: entity F port map(lamdaA => P(5)(847),lamdaB => P(5)(879),lamdaOut => P(4)(847));
U_F5848: entity F port map(lamdaA => P(5)(848),lamdaB => P(5)(880),lamdaOut => P(4)(848));
U_F5849: entity F port map(lamdaA => P(5)(849),lamdaB => P(5)(881),lamdaOut => P(4)(849));
U_F5850: entity F port map(lamdaA => P(5)(850),lamdaB => P(5)(882),lamdaOut => P(4)(850));
U_F5851: entity F port map(lamdaA => P(5)(851),lamdaB => P(5)(883),lamdaOut => P(4)(851));
U_F5852: entity F port map(lamdaA => P(5)(852),lamdaB => P(5)(884),lamdaOut => P(4)(852));
U_F5853: entity F port map(lamdaA => P(5)(853),lamdaB => P(5)(885),lamdaOut => P(4)(853));
U_F5854: entity F port map(lamdaA => P(5)(854),lamdaB => P(5)(886),lamdaOut => P(4)(854));
U_F5855: entity F port map(lamdaA => P(5)(855),lamdaB => P(5)(887),lamdaOut => P(4)(855));
U_F5856: entity F port map(lamdaA => P(5)(856),lamdaB => P(5)(888),lamdaOut => P(4)(856));
U_F5857: entity F port map(lamdaA => P(5)(857),lamdaB => P(5)(889),lamdaOut => P(4)(857));
U_F5858: entity F port map(lamdaA => P(5)(858),lamdaB => P(5)(890),lamdaOut => P(4)(858));
U_F5859: entity F port map(lamdaA => P(5)(859),lamdaB => P(5)(891),lamdaOut => P(4)(859));
U_F5860: entity F port map(lamdaA => P(5)(860),lamdaB => P(5)(892),lamdaOut => P(4)(860));
U_F5861: entity F port map(lamdaA => P(5)(861),lamdaB => P(5)(893),lamdaOut => P(4)(861));
U_F5862: entity F port map(lamdaA => P(5)(862),lamdaB => P(5)(894),lamdaOut => P(4)(862));
U_F5863: entity F port map(lamdaA => P(5)(863),lamdaB => P(5)(895),lamdaOut => P(4)(863));
U_G5864: entity G port map(lamdaA => P(5)(832),lamdaB => P(5)(864),s => s(5)(416),lamdaOut => P(4)(864));
U_G5865: entity G port map(lamdaA => P(5)(833),lamdaB => P(5)(865),s => s(5)(417),lamdaOut => P(4)(865));
U_G5866: entity G port map(lamdaA => P(5)(834),lamdaB => P(5)(866),s => s(5)(418),lamdaOut => P(4)(866));
U_G5867: entity G port map(lamdaA => P(5)(835),lamdaB => P(5)(867),s => s(5)(419),lamdaOut => P(4)(867));
U_G5868: entity G port map(lamdaA => P(5)(836),lamdaB => P(5)(868),s => s(5)(420),lamdaOut => P(4)(868));
U_G5869: entity G port map(lamdaA => P(5)(837),lamdaB => P(5)(869),s => s(5)(421),lamdaOut => P(4)(869));
U_G5870: entity G port map(lamdaA => P(5)(838),lamdaB => P(5)(870),s => s(5)(422),lamdaOut => P(4)(870));
U_G5871: entity G port map(lamdaA => P(5)(839),lamdaB => P(5)(871),s => s(5)(423),lamdaOut => P(4)(871));
U_G5872: entity G port map(lamdaA => P(5)(840),lamdaB => P(5)(872),s => s(5)(424),lamdaOut => P(4)(872));
U_G5873: entity G port map(lamdaA => P(5)(841),lamdaB => P(5)(873),s => s(5)(425),lamdaOut => P(4)(873));
U_G5874: entity G port map(lamdaA => P(5)(842),lamdaB => P(5)(874),s => s(5)(426),lamdaOut => P(4)(874));
U_G5875: entity G port map(lamdaA => P(5)(843),lamdaB => P(5)(875),s => s(5)(427),lamdaOut => P(4)(875));
U_G5876: entity G port map(lamdaA => P(5)(844),lamdaB => P(5)(876),s => s(5)(428),lamdaOut => P(4)(876));
U_G5877: entity G port map(lamdaA => P(5)(845),lamdaB => P(5)(877),s => s(5)(429),lamdaOut => P(4)(877));
U_G5878: entity G port map(lamdaA => P(5)(846),lamdaB => P(5)(878),s => s(5)(430),lamdaOut => P(4)(878));
U_G5879: entity G port map(lamdaA => P(5)(847),lamdaB => P(5)(879),s => s(5)(431),lamdaOut => P(4)(879));
U_G5880: entity G port map(lamdaA => P(5)(848),lamdaB => P(5)(880),s => s(5)(432),lamdaOut => P(4)(880));
U_G5881: entity G port map(lamdaA => P(5)(849),lamdaB => P(5)(881),s => s(5)(433),lamdaOut => P(4)(881));
U_G5882: entity G port map(lamdaA => P(5)(850),lamdaB => P(5)(882),s => s(5)(434),lamdaOut => P(4)(882));
U_G5883: entity G port map(lamdaA => P(5)(851),lamdaB => P(5)(883),s => s(5)(435),lamdaOut => P(4)(883));
U_G5884: entity G port map(lamdaA => P(5)(852),lamdaB => P(5)(884),s => s(5)(436),lamdaOut => P(4)(884));
U_G5885: entity G port map(lamdaA => P(5)(853),lamdaB => P(5)(885),s => s(5)(437),lamdaOut => P(4)(885));
U_G5886: entity G port map(lamdaA => P(5)(854),lamdaB => P(5)(886),s => s(5)(438),lamdaOut => P(4)(886));
U_G5887: entity G port map(lamdaA => P(5)(855),lamdaB => P(5)(887),s => s(5)(439),lamdaOut => P(4)(887));
U_G5888: entity G port map(lamdaA => P(5)(856),lamdaB => P(5)(888),s => s(5)(440),lamdaOut => P(4)(888));
U_G5889: entity G port map(lamdaA => P(5)(857),lamdaB => P(5)(889),s => s(5)(441),lamdaOut => P(4)(889));
U_G5890: entity G port map(lamdaA => P(5)(858),lamdaB => P(5)(890),s => s(5)(442),lamdaOut => P(4)(890));
U_G5891: entity G port map(lamdaA => P(5)(859),lamdaB => P(5)(891),s => s(5)(443),lamdaOut => P(4)(891));
U_G5892: entity G port map(lamdaA => P(5)(860),lamdaB => P(5)(892),s => s(5)(444),lamdaOut => P(4)(892));
U_G5893: entity G port map(lamdaA => P(5)(861),lamdaB => P(5)(893),s => s(5)(445),lamdaOut => P(4)(893));
U_G5894: entity G port map(lamdaA => P(5)(862),lamdaB => P(5)(894),s => s(5)(446),lamdaOut => P(4)(894));
U_G5895: entity G port map(lamdaA => P(5)(863),lamdaB => P(5)(895),s => s(5)(447),lamdaOut => P(4)(895));
U_F5896: entity F port map(lamdaA => P(5)(896),lamdaB => P(5)(928),lamdaOut => P(4)(896));
U_F5897: entity F port map(lamdaA => P(5)(897),lamdaB => P(5)(929),lamdaOut => P(4)(897));
U_F5898: entity F port map(lamdaA => P(5)(898),lamdaB => P(5)(930),lamdaOut => P(4)(898));
U_F5899: entity F port map(lamdaA => P(5)(899),lamdaB => P(5)(931),lamdaOut => P(4)(899));
U_F5900: entity F port map(lamdaA => P(5)(900),lamdaB => P(5)(932),lamdaOut => P(4)(900));
U_F5901: entity F port map(lamdaA => P(5)(901),lamdaB => P(5)(933),lamdaOut => P(4)(901));
U_F5902: entity F port map(lamdaA => P(5)(902),lamdaB => P(5)(934),lamdaOut => P(4)(902));
U_F5903: entity F port map(lamdaA => P(5)(903),lamdaB => P(5)(935),lamdaOut => P(4)(903));
U_F5904: entity F port map(lamdaA => P(5)(904),lamdaB => P(5)(936),lamdaOut => P(4)(904));
U_F5905: entity F port map(lamdaA => P(5)(905),lamdaB => P(5)(937),lamdaOut => P(4)(905));
U_F5906: entity F port map(lamdaA => P(5)(906),lamdaB => P(5)(938),lamdaOut => P(4)(906));
U_F5907: entity F port map(lamdaA => P(5)(907),lamdaB => P(5)(939),lamdaOut => P(4)(907));
U_F5908: entity F port map(lamdaA => P(5)(908),lamdaB => P(5)(940),lamdaOut => P(4)(908));
U_F5909: entity F port map(lamdaA => P(5)(909),lamdaB => P(5)(941),lamdaOut => P(4)(909));
U_F5910: entity F port map(lamdaA => P(5)(910),lamdaB => P(5)(942),lamdaOut => P(4)(910));
U_F5911: entity F port map(lamdaA => P(5)(911),lamdaB => P(5)(943),lamdaOut => P(4)(911));
U_F5912: entity F port map(lamdaA => P(5)(912),lamdaB => P(5)(944),lamdaOut => P(4)(912));
U_F5913: entity F port map(lamdaA => P(5)(913),lamdaB => P(5)(945),lamdaOut => P(4)(913));
U_F5914: entity F port map(lamdaA => P(5)(914),lamdaB => P(5)(946),lamdaOut => P(4)(914));
U_F5915: entity F port map(lamdaA => P(5)(915),lamdaB => P(5)(947),lamdaOut => P(4)(915));
U_F5916: entity F port map(lamdaA => P(5)(916),lamdaB => P(5)(948),lamdaOut => P(4)(916));
U_F5917: entity F port map(lamdaA => P(5)(917),lamdaB => P(5)(949),lamdaOut => P(4)(917));
U_F5918: entity F port map(lamdaA => P(5)(918),lamdaB => P(5)(950),lamdaOut => P(4)(918));
U_F5919: entity F port map(lamdaA => P(5)(919),lamdaB => P(5)(951),lamdaOut => P(4)(919));
U_F5920: entity F port map(lamdaA => P(5)(920),lamdaB => P(5)(952),lamdaOut => P(4)(920));
U_F5921: entity F port map(lamdaA => P(5)(921),lamdaB => P(5)(953),lamdaOut => P(4)(921));
U_F5922: entity F port map(lamdaA => P(5)(922),lamdaB => P(5)(954),lamdaOut => P(4)(922));
U_F5923: entity F port map(lamdaA => P(5)(923),lamdaB => P(5)(955),lamdaOut => P(4)(923));
U_F5924: entity F port map(lamdaA => P(5)(924),lamdaB => P(5)(956),lamdaOut => P(4)(924));
U_F5925: entity F port map(lamdaA => P(5)(925),lamdaB => P(5)(957),lamdaOut => P(4)(925));
U_F5926: entity F port map(lamdaA => P(5)(926),lamdaB => P(5)(958),lamdaOut => P(4)(926));
U_F5927: entity F port map(lamdaA => P(5)(927),lamdaB => P(5)(959),lamdaOut => P(4)(927));
U_G5928: entity G port map(lamdaA => P(5)(896),lamdaB => P(5)(928),s => s(5)(448),lamdaOut => P(4)(928));
U_G5929: entity G port map(lamdaA => P(5)(897),lamdaB => P(5)(929),s => s(5)(449),lamdaOut => P(4)(929));
U_G5930: entity G port map(lamdaA => P(5)(898),lamdaB => P(5)(930),s => s(5)(450),lamdaOut => P(4)(930));
U_G5931: entity G port map(lamdaA => P(5)(899),lamdaB => P(5)(931),s => s(5)(451),lamdaOut => P(4)(931));
U_G5932: entity G port map(lamdaA => P(5)(900),lamdaB => P(5)(932),s => s(5)(452),lamdaOut => P(4)(932));
U_G5933: entity G port map(lamdaA => P(5)(901),lamdaB => P(5)(933),s => s(5)(453),lamdaOut => P(4)(933));
U_G5934: entity G port map(lamdaA => P(5)(902),lamdaB => P(5)(934),s => s(5)(454),lamdaOut => P(4)(934));
U_G5935: entity G port map(lamdaA => P(5)(903),lamdaB => P(5)(935),s => s(5)(455),lamdaOut => P(4)(935));
U_G5936: entity G port map(lamdaA => P(5)(904),lamdaB => P(5)(936),s => s(5)(456),lamdaOut => P(4)(936));
U_G5937: entity G port map(lamdaA => P(5)(905),lamdaB => P(5)(937),s => s(5)(457),lamdaOut => P(4)(937));
U_G5938: entity G port map(lamdaA => P(5)(906),lamdaB => P(5)(938),s => s(5)(458),lamdaOut => P(4)(938));
U_G5939: entity G port map(lamdaA => P(5)(907),lamdaB => P(5)(939),s => s(5)(459),lamdaOut => P(4)(939));
U_G5940: entity G port map(lamdaA => P(5)(908),lamdaB => P(5)(940),s => s(5)(460),lamdaOut => P(4)(940));
U_G5941: entity G port map(lamdaA => P(5)(909),lamdaB => P(5)(941),s => s(5)(461),lamdaOut => P(4)(941));
U_G5942: entity G port map(lamdaA => P(5)(910),lamdaB => P(5)(942),s => s(5)(462),lamdaOut => P(4)(942));
U_G5943: entity G port map(lamdaA => P(5)(911),lamdaB => P(5)(943),s => s(5)(463),lamdaOut => P(4)(943));
U_G5944: entity G port map(lamdaA => P(5)(912),lamdaB => P(5)(944),s => s(5)(464),lamdaOut => P(4)(944));
U_G5945: entity G port map(lamdaA => P(5)(913),lamdaB => P(5)(945),s => s(5)(465),lamdaOut => P(4)(945));
U_G5946: entity G port map(lamdaA => P(5)(914),lamdaB => P(5)(946),s => s(5)(466),lamdaOut => P(4)(946));
U_G5947: entity G port map(lamdaA => P(5)(915),lamdaB => P(5)(947),s => s(5)(467),lamdaOut => P(4)(947));
U_G5948: entity G port map(lamdaA => P(5)(916),lamdaB => P(5)(948),s => s(5)(468),lamdaOut => P(4)(948));
U_G5949: entity G port map(lamdaA => P(5)(917),lamdaB => P(5)(949),s => s(5)(469),lamdaOut => P(4)(949));
U_G5950: entity G port map(lamdaA => P(5)(918),lamdaB => P(5)(950),s => s(5)(470),lamdaOut => P(4)(950));
U_G5951: entity G port map(lamdaA => P(5)(919),lamdaB => P(5)(951),s => s(5)(471),lamdaOut => P(4)(951));
U_G5952: entity G port map(lamdaA => P(5)(920),lamdaB => P(5)(952),s => s(5)(472),lamdaOut => P(4)(952));
U_G5953: entity G port map(lamdaA => P(5)(921),lamdaB => P(5)(953),s => s(5)(473),lamdaOut => P(4)(953));
U_G5954: entity G port map(lamdaA => P(5)(922),lamdaB => P(5)(954),s => s(5)(474),lamdaOut => P(4)(954));
U_G5955: entity G port map(lamdaA => P(5)(923),lamdaB => P(5)(955),s => s(5)(475),lamdaOut => P(4)(955));
U_G5956: entity G port map(lamdaA => P(5)(924),lamdaB => P(5)(956),s => s(5)(476),lamdaOut => P(4)(956));
U_G5957: entity G port map(lamdaA => P(5)(925),lamdaB => P(5)(957),s => s(5)(477),lamdaOut => P(4)(957));
U_G5958: entity G port map(lamdaA => P(5)(926),lamdaB => P(5)(958),s => s(5)(478),lamdaOut => P(4)(958));
U_G5959: entity G port map(lamdaA => P(5)(927),lamdaB => P(5)(959),s => s(5)(479),lamdaOut => P(4)(959));
U_F5960: entity F port map(lamdaA => P(5)(960),lamdaB => P(5)(992),lamdaOut => P(4)(960));
U_F5961: entity F port map(lamdaA => P(5)(961),lamdaB => P(5)(993),lamdaOut => P(4)(961));
U_F5962: entity F port map(lamdaA => P(5)(962),lamdaB => P(5)(994),lamdaOut => P(4)(962));
U_F5963: entity F port map(lamdaA => P(5)(963),lamdaB => P(5)(995),lamdaOut => P(4)(963));
U_F5964: entity F port map(lamdaA => P(5)(964),lamdaB => P(5)(996),lamdaOut => P(4)(964));
U_F5965: entity F port map(lamdaA => P(5)(965),lamdaB => P(5)(997),lamdaOut => P(4)(965));
U_F5966: entity F port map(lamdaA => P(5)(966),lamdaB => P(5)(998),lamdaOut => P(4)(966));
U_F5967: entity F port map(lamdaA => P(5)(967),lamdaB => P(5)(999),lamdaOut => P(4)(967));
U_F5968: entity F port map(lamdaA => P(5)(968),lamdaB => P(5)(1000),lamdaOut => P(4)(968));
U_F5969: entity F port map(lamdaA => P(5)(969),lamdaB => P(5)(1001),lamdaOut => P(4)(969));
U_F5970: entity F port map(lamdaA => P(5)(970),lamdaB => P(5)(1002),lamdaOut => P(4)(970));
U_F5971: entity F port map(lamdaA => P(5)(971),lamdaB => P(5)(1003),lamdaOut => P(4)(971));
U_F5972: entity F port map(lamdaA => P(5)(972),lamdaB => P(5)(1004),lamdaOut => P(4)(972));
U_F5973: entity F port map(lamdaA => P(5)(973),lamdaB => P(5)(1005),lamdaOut => P(4)(973));
U_F5974: entity F port map(lamdaA => P(5)(974),lamdaB => P(5)(1006),lamdaOut => P(4)(974));
U_F5975: entity F port map(lamdaA => P(5)(975),lamdaB => P(5)(1007),lamdaOut => P(4)(975));
U_F5976: entity F port map(lamdaA => P(5)(976),lamdaB => P(5)(1008),lamdaOut => P(4)(976));
U_F5977: entity F port map(lamdaA => P(5)(977),lamdaB => P(5)(1009),lamdaOut => P(4)(977));
U_F5978: entity F port map(lamdaA => P(5)(978),lamdaB => P(5)(1010),lamdaOut => P(4)(978));
U_F5979: entity F port map(lamdaA => P(5)(979),lamdaB => P(5)(1011),lamdaOut => P(4)(979));
U_F5980: entity F port map(lamdaA => P(5)(980),lamdaB => P(5)(1012),lamdaOut => P(4)(980));
U_F5981: entity F port map(lamdaA => P(5)(981),lamdaB => P(5)(1013),lamdaOut => P(4)(981));
U_F5982: entity F port map(lamdaA => P(5)(982),lamdaB => P(5)(1014),lamdaOut => P(4)(982));
U_F5983: entity F port map(lamdaA => P(5)(983),lamdaB => P(5)(1015),lamdaOut => P(4)(983));
U_F5984: entity F port map(lamdaA => P(5)(984),lamdaB => P(5)(1016),lamdaOut => P(4)(984));
U_F5985: entity F port map(lamdaA => P(5)(985),lamdaB => P(5)(1017),lamdaOut => P(4)(985));
U_F5986: entity F port map(lamdaA => P(5)(986),lamdaB => P(5)(1018),lamdaOut => P(4)(986));
U_F5987: entity F port map(lamdaA => P(5)(987),lamdaB => P(5)(1019),lamdaOut => P(4)(987));
U_F5988: entity F port map(lamdaA => P(5)(988),lamdaB => P(5)(1020),lamdaOut => P(4)(988));
U_F5989: entity F port map(lamdaA => P(5)(989),lamdaB => P(5)(1021),lamdaOut => P(4)(989));
U_F5990: entity F port map(lamdaA => P(5)(990),lamdaB => P(5)(1022),lamdaOut => P(4)(990));
U_F5991: entity F port map(lamdaA => P(5)(991),lamdaB => P(5)(1023),lamdaOut => P(4)(991));
U_G5992: entity G port map(lamdaA => P(5)(960),lamdaB => P(5)(992),s => s(5)(480),lamdaOut => P(4)(992));
U_G5993: entity G port map(lamdaA => P(5)(961),lamdaB => P(5)(993),s => s(5)(481),lamdaOut => P(4)(993));
U_G5994: entity G port map(lamdaA => P(5)(962),lamdaB => P(5)(994),s => s(5)(482),lamdaOut => P(4)(994));
U_G5995: entity G port map(lamdaA => P(5)(963),lamdaB => P(5)(995),s => s(5)(483),lamdaOut => P(4)(995));
U_G5996: entity G port map(lamdaA => P(5)(964),lamdaB => P(5)(996),s => s(5)(484),lamdaOut => P(4)(996));
U_G5997: entity G port map(lamdaA => P(5)(965),lamdaB => P(5)(997),s => s(5)(485),lamdaOut => P(4)(997));
U_G5998: entity G port map(lamdaA => P(5)(966),lamdaB => P(5)(998),s => s(5)(486),lamdaOut => P(4)(998));
U_G5999: entity G port map(lamdaA => P(5)(967),lamdaB => P(5)(999),s => s(5)(487),lamdaOut => P(4)(999));
U_G51000: entity G port map(lamdaA => P(5)(968),lamdaB => P(5)(1000),s => s(5)(488),lamdaOut => P(4)(1000));
U_G51001: entity G port map(lamdaA => P(5)(969),lamdaB => P(5)(1001),s => s(5)(489),lamdaOut => P(4)(1001));
U_G51002: entity G port map(lamdaA => P(5)(970),lamdaB => P(5)(1002),s => s(5)(490),lamdaOut => P(4)(1002));
U_G51003: entity G port map(lamdaA => P(5)(971),lamdaB => P(5)(1003),s => s(5)(491),lamdaOut => P(4)(1003));
U_G51004: entity G port map(lamdaA => P(5)(972),lamdaB => P(5)(1004),s => s(5)(492),lamdaOut => P(4)(1004));
U_G51005: entity G port map(lamdaA => P(5)(973),lamdaB => P(5)(1005),s => s(5)(493),lamdaOut => P(4)(1005));
U_G51006: entity G port map(lamdaA => P(5)(974),lamdaB => P(5)(1006),s => s(5)(494),lamdaOut => P(4)(1006));
U_G51007: entity G port map(lamdaA => P(5)(975),lamdaB => P(5)(1007),s => s(5)(495),lamdaOut => P(4)(1007));
U_G51008: entity G port map(lamdaA => P(5)(976),lamdaB => P(5)(1008),s => s(5)(496),lamdaOut => P(4)(1008));
U_G51009: entity G port map(lamdaA => P(5)(977),lamdaB => P(5)(1009),s => s(5)(497),lamdaOut => P(4)(1009));
U_G51010: entity G port map(lamdaA => P(5)(978),lamdaB => P(5)(1010),s => s(5)(498),lamdaOut => P(4)(1010));
U_G51011: entity G port map(lamdaA => P(5)(979),lamdaB => P(5)(1011),s => s(5)(499),lamdaOut => P(4)(1011));
U_G51012: entity G port map(lamdaA => P(5)(980),lamdaB => P(5)(1012),s => s(5)(500),lamdaOut => P(4)(1012));
U_G51013: entity G port map(lamdaA => P(5)(981),lamdaB => P(5)(1013),s => s(5)(501),lamdaOut => P(4)(1013));
U_G51014: entity G port map(lamdaA => P(5)(982),lamdaB => P(5)(1014),s => s(5)(502),lamdaOut => P(4)(1014));
U_G51015: entity G port map(lamdaA => P(5)(983),lamdaB => P(5)(1015),s => s(5)(503),lamdaOut => P(4)(1015));
U_G51016: entity G port map(lamdaA => P(5)(984),lamdaB => P(5)(1016),s => s(5)(504),lamdaOut => P(4)(1016));
U_G51017: entity G port map(lamdaA => P(5)(985),lamdaB => P(5)(1017),s => s(5)(505),lamdaOut => P(4)(1017));
U_G51018: entity G port map(lamdaA => P(5)(986),lamdaB => P(5)(1018),s => s(5)(506),lamdaOut => P(4)(1018));
U_G51019: entity G port map(lamdaA => P(5)(987),lamdaB => P(5)(1019),s => s(5)(507),lamdaOut => P(4)(1019));
U_G51020: entity G port map(lamdaA => P(5)(988),lamdaB => P(5)(1020),s => s(5)(508),lamdaOut => P(4)(1020));
U_G51021: entity G port map(lamdaA => P(5)(989),lamdaB => P(5)(1021),s => s(5)(509),lamdaOut => P(4)(1021));
U_G51022: entity G port map(lamdaA => P(5)(990),lamdaB => P(5)(1022),s => s(5)(510),lamdaOut => P(4)(1022));
U_G51023: entity G port map(lamdaA => P(5)(991),lamdaB => P(5)(1023),s => s(5)(511),lamdaOut => P(4)(1023));
-- STAGE 3
U_F40: entity F port map(lamdaA => P(4)(0),lamdaB => P(4)(64),lamdaOut => P(3)(0));
U_F41: entity F port map(lamdaA => P(4)(1),lamdaB => P(4)(65),lamdaOut => P(3)(1));
U_F42: entity F port map(lamdaA => P(4)(2),lamdaB => P(4)(66),lamdaOut => P(3)(2));
U_F43: entity F port map(lamdaA => P(4)(3),lamdaB => P(4)(67),lamdaOut => P(3)(3));
U_F44: entity F port map(lamdaA => P(4)(4),lamdaB => P(4)(68),lamdaOut => P(3)(4));
U_F45: entity F port map(lamdaA => P(4)(5),lamdaB => P(4)(69),lamdaOut => P(3)(5));
U_F46: entity F port map(lamdaA => P(4)(6),lamdaB => P(4)(70),lamdaOut => P(3)(6));
U_F47: entity F port map(lamdaA => P(4)(7),lamdaB => P(4)(71),lamdaOut => P(3)(7));
U_F48: entity F port map(lamdaA => P(4)(8),lamdaB => P(4)(72),lamdaOut => P(3)(8));
U_F49: entity F port map(lamdaA => P(4)(9),lamdaB => P(4)(73),lamdaOut => P(3)(9));
U_F410: entity F port map(lamdaA => P(4)(10),lamdaB => P(4)(74),lamdaOut => P(3)(10));
U_F411: entity F port map(lamdaA => P(4)(11),lamdaB => P(4)(75),lamdaOut => P(3)(11));
U_F412: entity F port map(lamdaA => P(4)(12),lamdaB => P(4)(76),lamdaOut => P(3)(12));
U_F413: entity F port map(lamdaA => P(4)(13),lamdaB => P(4)(77),lamdaOut => P(3)(13));
U_F414: entity F port map(lamdaA => P(4)(14),lamdaB => P(4)(78),lamdaOut => P(3)(14));
U_F415: entity F port map(lamdaA => P(4)(15),lamdaB => P(4)(79),lamdaOut => P(3)(15));
U_F416: entity F port map(lamdaA => P(4)(16),lamdaB => P(4)(80),lamdaOut => P(3)(16));
U_F417: entity F port map(lamdaA => P(4)(17),lamdaB => P(4)(81),lamdaOut => P(3)(17));
U_F418: entity F port map(lamdaA => P(4)(18),lamdaB => P(4)(82),lamdaOut => P(3)(18));
U_F419: entity F port map(lamdaA => P(4)(19),lamdaB => P(4)(83),lamdaOut => P(3)(19));
U_F420: entity F port map(lamdaA => P(4)(20),lamdaB => P(4)(84),lamdaOut => P(3)(20));
U_F421: entity F port map(lamdaA => P(4)(21),lamdaB => P(4)(85),lamdaOut => P(3)(21));
U_F422: entity F port map(lamdaA => P(4)(22),lamdaB => P(4)(86),lamdaOut => P(3)(22));
U_F423: entity F port map(lamdaA => P(4)(23),lamdaB => P(4)(87),lamdaOut => P(3)(23));
U_F424: entity F port map(lamdaA => P(4)(24),lamdaB => P(4)(88),lamdaOut => P(3)(24));
U_F425: entity F port map(lamdaA => P(4)(25),lamdaB => P(4)(89),lamdaOut => P(3)(25));
U_F426: entity F port map(lamdaA => P(4)(26),lamdaB => P(4)(90),lamdaOut => P(3)(26));
U_F427: entity F port map(lamdaA => P(4)(27),lamdaB => P(4)(91),lamdaOut => P(3)(27));
U_F428: entity F port map(lamdaA => P(4)(28),lamdaB => P(4)(92),lamdaOut => P(3)(28));
U_F429: entity F port map(lamdaA => P(4)(29),lamdaB => P(4)(93),lamdaOut => P(3)(29));
U_F430: entity F port map(lamdaA => P(4)(30),lamdaB => P(4)(94),lamdaOut => P(3)(30));
U_F431: entity F port map(lamdaA => P(4)(31),lamdaB => P(4)(95),lamdaOut => P(3)(31));
U_F432: entity F port map(lamdaA => P(4)(32),lamdaB => P(4)(96),lamdaOut => P(3)(32));
U_F433: entity F port map(lamdaA => P(4)(33),lamdaB => P(4)(97),lamdaOut => P(3)(33));
U_F434: entity F port map(lamdaA => P(4)(34),lamdaB => P(4)(98),lamdaOut => P(3)(34));
U_F435: entity F port map(lamdaA => P(4)(35),lamdaB => P(4)(99),lamdaOut => P(3)(35));
U_F436: entity F port map(lamdaA => P(4)(36),lamdaB => P(4)(100),lamdaOut => P(3)(36));
U_F437: entity F port map(lamdaA => P(4)(37),lamdaB => P(4)(101),lamdaOut => P(3)(37));
U_F438: entity F port map(lamdaA => P(4)(38),lamdaB => P(4)(102),lamdaOut => P(3)(38));
U_F439: entity F port map(lamdaA => P(4)(39),lamdaB => P(4)(103),lamdaOut => P(3)(39));
U_F440: entity F port map(lamdaA => P(4)(40),lamdaB => P(4)(104),lamdaOut => P(3)(40));
U_F441: entity F port map(lamdaA => P(4)(41),lamdaB => P(4)(105),lamdaOut => P(3)(41));
U_F442: entity F port map(lamdaA => P(4)(42),lamdaB => P(4)(106),lamdaOut => P(3)(42));
U_F443: entity F port map(lamdaA => P(4)(43),lamdaB => P(4)(107),lamdaOut => P(3)(43));
U_F444: entity F port map(lamdaA => P(4)(44),lamdaB => P(4)(108),lamdaOut => P(3)(44));
U_F445: entity F port map(lamdaA => P(4)(45),lamdaB => P(4)(109),lamdaOut => P(3)(45));
U_F446: entity F port map(lamdaA => P(4)(46),lamdaB => P(4)(110),lamdaOut => P(3)(46));
U_F447: entity F port map(lamdaA => P(4)(47),lamdaB => P(4)(111),lamdaOut => P(3)(47));
U_F448: entity F port map(lamdaA => P(4)(48),lamdaB => P(4)(112),lamdaOut => P(3)(48));
U_F449: entity F port map(lamdaA => P(4)(49),lamdaB => P(4)(113),lamdaOut => P(3)(49));
U_F450: entity F port map(lamdaA => P(4)(50),lamdaB => P(4)(114),lamdaOut => P(3)(50));
U_F451: entity F port map(lamdaA => P(4)(51),lamdaB => P(4)(115),lamdaOut => P(3)(51));
U_F452: entity F port map(lamdaA => P(4)(52),lamdaB => P(4)(116),lamdaOut => P(3)(52));
U_F453: entity F port map(lamdaA => P(4)(53),lamdaB => P(4)(117),lamdaOut => P(3)(53));
U_F454: entity F port map(lamdaA => P(4)(54),lamdaB => P(4)(118),lamdaOut => P(3)(54));
U_F455: entity F port map(lamdaA => P(4)(55),lamdaB => P(4)(119),lamdaOut => P(3)(55));
U_F456: entity F port map(lamdaA => P(4)(56),lamdaB => P(4)(120),lamdaOut => P(3)(56));
U_F457: entity F port map(lamdaA => P(4)(57),lamdaB => P(4)(121),lamdaOut => P(3)(57));
U_F458: entity F port map(lamdaA => P(4)(58),lamdaB => P(4)(122),lamdaOut => P(3)(58));
U_F459: entity F port map(lamdaA => P(4)(59),lamdaB => P(4)(123),lamdaOut => P(3)(59));
U_F460: entity F port map(lamdaA => P(4)(60),lamdaB => P(4)(124),lamdaOut => P(3)(60));
U_F461: entity F port map(lamdaA => P(4)(61),lamdaB => P(4)(125),lamdaOut => P(3)(61));
U_F462: entity F port map(lamdaA => P(4)(62),lamdaB => P(4)(126),lamdaOut => P(3)(62));
U_F463: entity F port map(lamdaA => P(4)(63),lamdaB => P(4)(127),lamdaOut => P(3)(63));
U_G464: entity G port map(lamdaA => P(4)(0),lamdaB => P(4)(64),s => s(4)(0),lamdaOut => P(3)(64));
U_G465: entity G port map(lamdaA => P(4)(1),lamdaB => P(4)(65),s => s(4)(1),lamdaOut => P(3)(65));
U_G466: entity G port map(lamdaA => P(4)(2),lamdaB => P(4)(66),s => s(4)(2),lamdaOut => P(3)(66));
U_G467: entity G port map(lamdaA => P(4)(3),lamdaB => P(4)(67),s => s(4)(3),lamdaOut => P(3)(67));
U_G468: entity G port map(lamdaA => P(4)(4),lamdaB => P(4)(68),s => s(4)(4),lamdaOut => P(3)(68));
U_G469: entity G port map(lamdaA => P(4)(5),lamdaB => P(4)(69),s => s(4)(5),lamdaOut => P(3)(69));
U_G470: entity G port map(lamdaA => P(4)(6),lamdaB => P(4)(70),s => s(4)(6),lamdaOut => P(3)(70));
U_G471: entity G port map(lamdaA => P(4)(7),lamdaB => P(4)(71),s => s(4)(7),lamdaOut => P(3)(71));
U_G472: entity G port map(lamdaA => P(4)(8),lamdaB => P(4)(72),s => s(4)(8),lamdaOut => P(3)(72));
U_G473: entity G port map(lamdaA => P(4)(9),lamdaB => P(4)(73),s => s(4)(9),lamdaOut => P(3)(73));
U_G474: entity G port map(lamdaA => P(4)(10),lamdaB => P(4)(74),s => s(4)(10),lamdaOut => P(3)(74));
U_G475: entity G port map(lamdaA => P(4)(11),lamdaB => P(4)(75),s => s(4)(11),lamdaOut => P(3)(75));
U_G476: entity G port map(lamdaA => P(4)(12),lamdaB => P(4)(76),s => s(4)(12),lamdaOut => P(3)(76));
U_G477: entity G port map(lamdaA => P(4)(13),lamdaB => P(4)(77),s => s(4)(13),lamdaOut => P(3)(77));
U_G478: entity G port map(lamdaA => P(4)(14),lamdaB => P(4)(78),s => s(4)(14),lamdaOut => P(3)(78));
U_G479: entity G port map(lamdaA => P(4)(15),lamdaB => P(4)(79),s => s(4)(15),lamdaOut => P(3)(79));
U_G480: entity G port map(lamdaA => P(4)(16),lamdaB => P(4)(80),s => s(4)(16),lamdaOut => P(3)(80));
U_G481: entity G port map(lamdaA => P(4)(17),lamdaB => P(4)(81),s => s(4)(17),lamdaOut => P(3)(81));
U_G482: entity G port map(lamdaA => P(4)(18),lamdaB => P(4)(82),s => s(4)(18),lamdaOut => P(3)(82));
U_G483: entity G port map(lamdaA => P(4)(19),lamdaB => P(4)(83),s => s(4)(19),lamdaOut => P(3)(83));
U_G484: entity G port map(lamdaA => P(4)(20),lamdaB => P(4)(84),s => s(4)(20),lamdaOut => P(3)(84));
U_G485: entity G port map(lamdaA => P(4)(21),lamdaB => P(4)(85),s => s(4)(21),lamdaOut => P(3)(85));
U_G486: entity G port map(lamdaA => P(4)(22),lamdaB => P(4)(86),s => s(4)(22),lamdaOut => P(3)(86));
U_G487: entity G port map(lamdaA => P(4)(23),lamdaB => P(4)(87),s => s(4)(23),lamdaOut => P(3)(87));
U_G488: entity G port map(lamdaA => P(4)(24),lamdaB => P(4)(88),s => s(4)(24),lamdaOut => P(3)(88));
U_G489: entity G port map(lamdaA => P(4)(25),lamdaB => P(4)(89),s => s(4)(25),lamdaOut => P(3)(89));
U_G490: entity G port map(lamdaA => P(4)(26),lamdaB => P(4)(90),s => s(4)(26),lamdaOut => P(3)(90));
U_G491: entity G port map(lamdaA => P(4)(27),lamdaB => P(4)(91),s => s(4)(27),lamdaOut => P(3)(91));
U_G492: entity G port map(lamdaA => P(4)(28),lamdaB => P(4)(92),s => s(4)(28),lamdaOut => P(3)(92));
U_G493: entity G port map(lamdaA => P(4)(29),lamdaB => P(4)(93),s => s(4)(29),lamdaOut => P(3)(93));
U_G494: entity G port map(lamdaA => P(4)(30),lamdaB => P(4)(94),s => s(4)(30),lamdaOut => P(3)(94));
U_G495: entity G port map(lamdaA => P(4)(31),lamdaB => P(4)(95),s => s(4)(31),lamdaOut => P(3)(95));
U_G496: entity G port map(lamdaA => P(4)(32),lamdaB => P(4)(96),s => s(4)(32),lamdaOut => P(3)(96));
U_G497: entity G port map(lamdaA => P(4)(33),lamdaB => P(4)(97),s => s(4)(33),lamdaOut => P(3)(97));
U_G498: entity G port map(lamdaA => P(4)(34),lamdaB => P(4)(98),s => s(4)(34),lamdaOut => P(3)(98));
U_G499: entity G port map(lamdaA => P(4)(35),lamdaB => P(4)(99),s => s(4)(35),lamdaOut => P(3)(99));
U_G4100: entity G port map(lamdaA => P(4)(36),lamdaB => P(4)(100),s => s(4)(36),lamdaOut => P(3)(100));
U_G4101: entity G port map(lamdaA => P(4)(37),lamdaB => P(4)(101),s => s(4)(37),lamdaOut => P(3)(101));
U_G4102: entity G port map(lamdaA => P(4)(38),lamdaB => P(4)(102),s => s(4)(38),lamdaOut => P(3)(102));
U_G4103: entity G port map(lamdaA => P(4)(39),lamdaB => P(4)(103),s => s(4)(39),lamdaOut => P(3)(103));
U_G4104: entity G port map(lamdaA => P(4)(40),lamdaB => P(4)(104),s => s(4)(40),lamdaOut => P(3)(104));
U_G4105: entity G port map(lamdaA => P(4)(41),lamdaB => P(4)(105),s => s(4)(41),lamdaOut => P(3)(105));
U_G4106: entity G port map(lamdaA => P(4)(42),lamdaB => P(4)(106),s => s(4)(42),lamdaOut => P(3)(106));
U_G4107: entity G port map(lamdaA => P(4)(43),lamdaB => P(4)(107),s => s(4)(43),lamdaOut => P(3)(107));
U_G4108: entity G port map(lamdaA => P(4)(44),lamdaB => P(4)(108),s => s(4)(44),lamdaOut => P(3)(108));
U_G4109: entity G port map(lamdaA => P(4)(45),lamdaB => P(4)(109),s => s(4)(45),lamdaOut => P(3)(109));
U_G4110: entity G port map(lamdaA => P(4)(46),lamdaB => P(4)(110),s => s(4)(46),lamdaOut => P(3)(110));
U_G4111: entity G port map(lamdaA => P(4)(47),lamdaB => P(4)(111),s => s(4)(47),lamdaOut => P(3)(111));
U_G4112: entity G port map(lamdaA => P(4)(48),lamdaB => P(4)(112),s => s(4)(48),lamdaOut => P(3)(112));
U_G4113: entity G port map(lamdaA => P(4)(49),lamdaB => P(4)(113),s => s(4)(49),lamdaOut => P(3)(113));
U_G4114: entity G port map(lamdaA => P(4)(50),lamdaB => P(4)(114),s => s(4)(50),lamdaOut => P(3)(114));
U_G4115: entity G port map(lamdaA => P(4)(51),lamdaB => P(4)(115),s => s(4)(51),lamdaOut => P(3)(115));
U_G4116: entity G port map(lamdaA => P(4)(52),lamdaB => P(4)(116),s => s(4)(52),lamdaOut => P(3)(116));
U_G4117: entity G port map(lamdaA => P(4)(53),lamdaB => P(4)(117),s => s(4)(53),lamdaOut => P(3)(117));
U_G4118: entity G port map(lamdaA => P(4)(54),lamdaB => P(4)(118),s => s(4)(54),lamdaOut => P(3)(118));
U_G4119: entity G port map(lamdaA => P(4)(55),lamdaB => P(4)(119),s => s(4)(55),lamdaOut => P(3)(119));
U_G4120: entity G port map(lamdaA => P(4)(56),lamdaB => P(4)(120),s => s(4)(56),lamdaOut => P(3)(120));
U_G4121: entity G port map(lamdaA => P(4)(57),lamdaB => P(4)(121),s => s(4)(57),lamdaOut => P(3)(121));
U_G4122: entity G port map(lamdaA => P(4)(58),lamdaB => P(4)(122),s => s(4)(58),lamdaOut => P(3)(122));
U_G4123: entity G port map(lamdaA => P(4)(59),lamdaB => P(4)(123),s => s(4)(59),lamdaOut => P(3)(123));
U_G4124: entity G port map(lamdaA => P(4)(60),lamdaB => P(4)(124),s => s(4)(60),lamdaOut => P(3)(124));
U_G4125: entity G port map(lamdaA => P(4)(61),lamdaB => P(4)(125),s => s(4)(61),lamdaOut => P(3)(125));
U_G4126: entity G port map(lamdaA => P(4)(62),lamdaB => P(4)(126),s => s(4)(62),lamdaOut => P(3)(126));
U_G4127: entity G port map(lamdaA => P(4)(63),lamdaB => P(4)(127),s => s(4)(63),lamdaOut => P(3)(127));
U_F4128: entity F port map(lamdaA => P(4)(128),lamdaB => P(4)(192),lamdaOut => P(3)(128));
U_F4129: entity F port map(lamdaA => P(4)(129),lamdaB => P(4)(193),lamdaOut => P(3)(129));
U_F4130: entity F port map(lamdaA => P(4)(130),lamdaB => P(4)(194),lamdaOut => P(3)(130));
U_F4131: entity F port map(lamdaA => P(4)(131),lamdaB => P(4)(195),lamdaOut => P(3)(131));
U_F4132: entity F port map(lamdaA => P(4)(132),lamdaB => P(4)(196),lamdaOut => P(3)(132));
U_F4133: entity F port map(lamdaA => P(4)(133),lamdaB => P(4)(197),lamdaOut => P(3)(133));
U_F4134: entity F port map(lamdaA => P(4)(134),lamdaB => P(4)(198),lamdaOut => P(3)(134));
U_F4135: entity F port map(lamdaA => P(4)(135),lamdaB => P(4)(199),lamdaOut => P(3)(135));
U_F4136: entity F port map(lamdaA => P(4)(136),lamdaB => P(4)(200),lamdaOut => P(3)(136));
U_F4137: entity F port map(lamdaA => P(4)(137),lamdaB => P(4)(201),lamdaOut => P(3)(137));
U_F4138: entity F port map(lamdaA => P(4)(138),lamdaB => P(4)(202),lamdaOut => P(3)(138));
U_F4139: entity F port map(lamdaA => P(4)(139),lamdaB => P(4)(203),lamdaOut => P(3)(139));
U_F4140: entity F port map(lamdaA => P(4)(140),lamdaB => P(4)(204),lamdaOut => P(3)(140));
U_F4141: entity F port map(lamdaA => P(4)(141),lamdaB => P(4)(205),lamdaOut => P(3)(141));
U_F4142: entity F port map(lamdaA => P(4)(142),lamdaB => P(4)(206),lamdaOut => P(3)(142));
U_F4143: entity F port map(lamdaA => P(4)(143),lamdaB => P(4)(207),lamdaOut => P(3)(143));
U_F4144: entity F port map(lamdaA => P(4)(144),lamdaB => P(4)(208),lamdaOut => P(3)(144));
U_F4145: entity F port map(lamdaA => P(4)(145),lamdaB => P(4)(209),lamdaOut => P(3)(145));
U_F4146: entity F port map(lamdaA => P(4)(146),lamdaB => P(4)(210),lamdaOut => P(3)(146));
U_F4147: entity F port map(lamdaA => P(4)(147),lamdaB => P(4)(211),lamdaOut => P(3)(147));
U_F4148: entity F port map(lamdaA => P(4)(148),lamdaB => P(4)(212),lamdaOut => P(3)(148));
U_F4149: entity F port map(lamdaA => P(4)(149),lamdaB => P(4)(213),lamdaOut => P(3)(149));
U_F4150: entity F port map(lamdaA => P(4)(150),lamdaB => P(4)(214),lamdaOut => P(3)(150));
U_F4151: entity F port map(lamdaA => P(4)(151),lamdaB => P(4)(215),lamdaOut => P(3)(151));
U_F4152: entity F port map(lamdaA => P(4)(152),lamdaB => P(4)(216),lamdaOut => P(3)(152));
U_F4153: entity F port map(lamdaA => P(4)(153),lamdaB => P(4)(217),lamdaOut => P(3)(153));
U_F4154: entity F port map(lamdaA => P(4)(154),lamdaB => P(4)(218),lamdaOut => P(3)(154));
U_F4155: entity F port map(lamdaA => P(4)(155),lamdaB => P(4)(219),lamdaOut => P(3)(155));
U_F4156: entity F port map(lamdaA => P(4)(156),lamdaB => P(4)(220),lamdaOut => P(3)(156));
U_F4157: entity F port map(lamdaA => P(4)(157),lamdaB => P(4)(221),lamdaOut => P(3)(157));
U_F4158: entity F port map(lamdaA => P(4)(158),lamdaB => P(4)(222),lamdaOut => P(3)(158));
U_F4159: entity F port map(lamdaA => P(4)(159),lamdaB => P(4)(223),lamdaOut => P(3)(159));
U_F4160: entity F port map(lamdaA => P(4)(160),lamdaB => P(4)(224),lamdaOut => P(3)(160));
U_F4161: entity F port map(lamdaA => P(4)(161),lamdaB => P(4)(225),lamdaOut => P(3)(161));
U_F4162: entity F port map(lamdaA => P(4)(162),lamdaB => P(4)(226),lamdaOut => P(3)(162));
U_F4163: entity F port map(lamdaA => P(4)(163),lamdaB => P(4)(227),lamdaOut => P(3)(163));
U_F4164: entity F port map(lamdaA => P(4)(164),lamdaB => P(4)(228),lamdaOut => P(3)(164));
U_F4165: entity F port map(lamdaA => P(4)(165),lamdaB => P(4)(229),lamdaOut => P(3)(165));
U_F4166: entity F port map(lamdaA => P(4)(166),lamdaB => P(4)(230),lamdaOut => P(3)(166));
U_F4167: entity F port map(lamdaA => P(4)(167),lamdaB => P(4)(231),lamdaOut => P(3)(167));
U_F4168: entity F port map(lamdaA => P(4)(168),lamdaB => P(4)(232),lamdaOut => P(3)(168));
U_F4169: entity F port map(lamdaA => P(4)(169),lamdaB => P(4)(233),lamdaOut => P(3)(169));
U_F4170: entity F port map(lamdaA => P(4)(170),lamdaB => P(4)(234),lamdaOut => P(3)(170));
U_F4171: entity F port map(lamdaA => P(4)(171),lamdaB => P(4)(235),lamdaOut => P(3)(171));
U_F4172: entity F port map(lamdaA => P(4)(172),lamdaB => P(4)(236),lamdaOut => P(3)(172));
U_F4173: entity F port map(lamdaA => P(4)(173),lamdaB => P(4)(237),lamdaOut => P(3)(173));
U_F4174: entity F port map(lamdaA => P(4)(174),lamdaB => P(4)(238),lamdaOut => P(3)(174));
U_F4175: entity F port map(lamdaA => P(4)(175),lamdaB => P(4)(239),lamdaOut => P(3)(175));
U_F4176: entity F port map(lamdaA => P(4)(176),lamdaB => P(4)(240),lamdaOut => P(3)(176));
U_F4177: entity F port map(lamdaA => P(4)(177),lamdaB => P(4)(241),lamdaOut => P(3)(177));
U_F4178: entity F port map(lamdaA => P(4)(178),lamdaB => P(4)(242),lamdaOut => P(3)(178));
U_F4179: entity F port map(lamdaA => P(4)(179),lamdaB => P(4)(243),lamdaOut => P(3)(179));
U_F4180: entity F port map(lamdaA => P(4)(180),lamdaB => P(4)(244),lamdaOut => P(3)(180));
U_F4181: entity F port map(lamdaA => P(4)(181),lamdaB => P(4)(245),lamdaOut => P(3)(181));
U_F4182: entity F port map(lamdaA => P(4)(182),lamdaB => P(4)(246),lamdaOut => P(3)(182));
U_F4183: entity F port map(lamdaA => P(4)(183),lamdaB => P(4)(247),lamdaOut => P(3)(183));
U_F4184: entity F port map(lamdaA => P(4)(184),lamdaB => P(4)(248),lamdaOut => P(3)(184));
U_F4185: entity F port map(lamdaA => P(4)(185),lamdaB => P(4)(249),lamdaOut => P(3)(185));
U_F4186: entity F port map(lamdaA => P(4)(186),lamdaB => P(4)(250),lamdaOut => P(3)(186));
U_F4187: entity F port map(lamdaA => P(4)(187),lamdaB => P(4)(251),lamdaOut => P(3)(187));
U_F4188: entity F port map(lamdaA => P(4)(188),lamdaB => P(4)(252),lamdaOut => P(3)(188));
U_F4189: entity F port map(lamdaA => P(4)(189),lamdaB => P(4)(253),lamdaOut => P(3)(189));
U_F4190: entity F port map(lamdaA => P(4)(190),lamdaB => P(4)(254),lamdaOut => P(3)(190));
U_F4191: entity F port map(lamdaA => P(4)(191),lamdaB => P(4)(255),lamdaOut => P(3)(191));
U_G4192: entity G port map(lamdaA => P(4)(128),lamdaB => P(4)(192),s => s(4)(64),lamdaOut => P(3)(192));
U_G4193: entity G port map(lamdaA => P(4)(129),lamdaB => P(4)(193),s => s(4)(65),lamdaOut => P(3)(193));
U_G4194: entity G port map(lamdaA => P(4)(130),lamdaB => P(4)(194),s => s(4)(66),lamdaOut => P(3)(194));
U_G4195: entity G port map(lamdaA => P(4)(131),lamdaB => P(4)(195),s => s(4)(67),lamdaOut => P(3)(195));
U_G4196: entity G port map(lamdaA => P(4)(132),lamdaB => P(4)(196),s => s(4)(68),lamdaOut => P(3)(196));
U_G4197: entity G port map(lamdaA => P(4)(133),lamdaB => P(4)(197),s => s(4)(69),lamdaOut => P(3)(197));
U_G4198: entity G port map(lamdaA => P(4)(134),lamdaB => P(4)(198),s => s(4)(70),lamdaOut => P(3)(198));
U_G4199: entity G port map(lamdaA => P(4)(135),lamdaB => P(4)(199),s => s(4)(71),lamdaOut => P(3)(199));
U_G4200: entity G port map(lamdaA => P(4)(136),lamdaB => P(4)(200),s => s(4)(72),lamdaOut => P(3)(200));
U_G4201: entity G port map(lamdaA => P(4)(137),lamdaB => P(4)(201),s => s(4)(73),lamdaOut => P(3)(201));
U_G4202: entity G port map(lamdaA => P(4)(138),lamdaB => P(4)(202),s => s(4)(74),lamdaOut => P(3)(202));
U_G4203: entity G port map(lamdaA => P(4)(139),lamdaB => P(4)(203),s => s(4)(75),lamdaOut => P(3)(203));
U_G4204: entity G port map(lamdaA => P(4)(140),lamdaB => P(4)(204),s => s(4)(76),lamdaOut => P(3)(204));
U_G4205: entity G port map(lamdaA => P(4)(141),lamdaB => P(4)(205),s => s(4)(77),lamdaOut => P(3)(205));
U_G4206: entity G port map(lamdaA => P(4)(142),lamdaB => P(4)(206),s => s(4)(78),lamdaOut => P(3)(206));
U_G4207: entity G port map(lamdaA => P(4)(143),lamdaB => P(4)(207),s => s(4)(79),lamdaOut => P(3)(207));
U_G4208: entity G port map(lamdaA => P(4)(144),lamdaB => P(4)(208),s => s(4)(80),lamdaOut => P(3)(208));
U_G4209: entity G port map(lamdaA => P(4)(145),lamdaB => P(4)(209),s => s(4)(81),lamdaOut => P(3)(209));
U_G4210: entity G port map(lamdaA => P(4)(146),lamdaB => P(4)(210),s => s(4)(82),lamdaOut => P(3)(210));
U_G4211: entity G port map(lamdaA => P(4)(147),lamdaB => P(4)(211),s => s(4)(83),lamdaOut => P(3)(211));
U_G4212: entity G port map(lamdaA => P(4)(148),lamdaB => P(4)(212),s => s(4)(84),lamdaOut => P(3)(212));
U_G4213: entity G port map(lamdaA => P(4)(149),lamdaB => P(4)(213),s => s(4)(85),lamdaOut => P(3)(213));
U_G4214: entity G port map(lamdaA => P(4)(150),lamdaB => P(4)(214),s => s(4)(86),lamdaOut => P(3)(214));
U_G4215: entity G port map(lamdaA => P(4)(151),lamdaB => P(4)(215),s => s(4)(87),lamdaOut => P(3)(215));
U_G4216: entity G port map(lamdaA => P(4)(152),lamdaB => P(4)(216),s => s(4)(88),lamdaOut => P(3)(216));
U_G4217: entity G port map(lamdaA => P(4)(153),lamdaB => P(4)(217),s => s(4)(89),lamdaOut => P(3)(217));
U_G4218: entity G port map(lamdaA => P(4)(154),lamdaB => P(4)(218),s => s(4)(90),lamdaOut => P(3)(218));
U_G4219: entity G port map(lamdaA => P(4)(155),lamdaB => P(4)(219),s => s(4)(91),lamdaOut => P(3)(219));
U_G4220: entity G port map(lamdaA => P(4)(156),lamdaB => P(4)(220),s => s(4)(92),lamdaOut => P(3)(220));
U_G4221: entity G port map(lamdaA => P(4)(157),lamdaB => P(4)(221),s => s(4)(93),lamdaOut => P(3)(221));
U_G4222: entity G port map(lamdaA => P(4)(158),lamdaB => P(4)(222),s => s(4)(94),lamdaOut => P(3)(222));
U_G4223: entity G port map(lamdaA => P(4)(159),lamdaB => P(4)(223),s => s(4)(95),lamdaOut => P(3)(223));
U_G4224: entity G port map(lamdaA => P(4)(160),lamdaB => P(4)(224),s => s(4)(96),lamdaOut => P(3)(224));
U_G4225: entity G port map(lamdaA => P(4)(161),lamdaB => P(4)(225),s => s(4)(97),lamdaOut => P(3)(225));
U_G4226: entity G port map(lamdaA => P(4)(162),lamdaB => P(4)(226),s => s(4)(98),lamdaOut => P(3)(226));
U_G4227: entity G port map(lamdaA => P(4)(163),lamdaB => P(4)(227),s => s(4)(99),lamdaOut => P(3)(227));
U_G4228: entity G port map(lamdaA => P(4)(164),lamdaB => P(4)(228),s => s(4)(100),lamdaOut => P(3)(228));
U_G4229: entity G port map(lamdaA => P(4)(165),lamdaB => P(4)(229),s => s(4)(101),lamdaOut => P(3)(229));
U_G4230: entity G port map(lamdaA => P(4)(166),lamdaB => P(4)(230),s => s(4)(102),lamdaOut => P(3)(230));
U_G4231: entity G port map(lamdaA => P(4)(167),lamdaB => P(4)(231),s => s(4)(103),lamdaOut => P(3)(231));
U_G4232: entity G port map(lamdaA => P(4)(168),lamdaB => P(4)(232),s => s(4)(104),lamdaOut => P(3)(232));
U_G4233: entity G port map(lamdaA => P(4)(169),lamdaB => P(4)(233),s => s(4)(105),lamdaOut => P(3)(233));
U_G4234: entity G port map(lamdaA => P(4)(170),lamdaB => P(4)(234),s => s(4)(106),lamdaOut => P(3)(234));
U_G4235: entity G port map(lamdaA => P(4)(171),lamdaB => P(4)(235),s => s(4)(107),lamdaOut => P(3)(235));
U_G4236: entity G port map(lamdaA => P(4)(172),lamdaB => P(4)(236),s => s(4)(108),lamdaOut => P(3)(236));
U_G4237: entity G port map(lamdaA => P(4)(173),lamdaB => P(4)(237),s => s(4)(109),lamdaOut => P(3)(237));
U_G4238: entity G port map(lamdaA => P(4)(174),lamdaB => P(4)(238),s => s(4)(110),lamdaOut => P(3)(238));
U_G4239: entity G port map(lamdaA => P(4)(175),lamdaB => P(4)(239),s => s(4)(111),lamdaOut => P(3)(239));
U_G4240: entity G port map(lamdaA => P(4)(176),lamdaB => P(4)(240),s => s(4)(112),lamdaOut => P(3)(240));
U_G4241: entity G port map(lamdaA => P(4)(177),lamdaB => P(4)(241),s => s(4)(113),lamdaOut => P(3)(241));
U_G4242: entity G port map(lamdaA => P(4)(178),lamdaB => P(4)(242),s => s(4)(114),lamdaOut => P(3)(242));
U_G4243: entity G port map(lamdaA => P(4)(179),lamdaB => P(4)(243),s => s(4)(115),lamdaOut => P(3)(243));
U_G4244: entity G port map(lamdaA => P(4)(180),lamdaB => P(4)(244),s => s(4)(116),lamdaOut => P(3)(244));
U_G4245: entity G port map(lamdaA => P(4)(181),lamdaB => P(4)(245),s => s(4)(117),lamdaOut => P(3)(245));
U_G4246: entity G port map(lamdaA => P(4)(182),lamdaB => P(4)(246),s => s(4)(118),lamdaOut => P(3)(246));
U_G4247: entity G port map(lamdaA => P(4)(183),lamdaB => P(4)(247),s => s(4)(119),lamdaOut => P(3)(247));
U_G4248: entity G port map(lamdaA => P(4)(184),lamdaB => P(4)(248),s => s(4)(120),lamdaOut => P(3)(248));
U_G4249: entity G port map(lamdaA => P(4)(185),lamdaB => P(4)(249),s => s(4)(121),lamdaOut => P(3)(249));
U_G4250: entity G port map(lamdaA => P(4)(186),lamdaB => P(4)(250),s => s(4)(122),lamdaOut => P(3)(250));
U_G4251: entity G port map(lamdaA => P(4)(187),lamdaB => P(4)(251),s => s(4)(123),lamdaOut => P(3)(251));
U_G4252: entity G port map(lamdaA => P(4)(188),lamdaB => P(4)(252),s => s(4)(124),lamdaOut => P(3)(252));
U_G4253: entity G port map(lamdaA => P(4)(189),lamdaB => P(4)(253),s => s(4)(125),lamdaOut => P(3)(253));
U_G4254: entity G port map(lamdaA => P(4)(190),lamdaB => P(4)(254),s => s(4)(126),lamdaOut => P(3)(254));
U_G4255: entity G port map(lamdaA => P(4)(191),lamdaB => P(4)(255),s => s(4)(127),lamdaOut => P(3)(255));
U_F4256: entity F port map(lamdaA => P(4)(256),lamdaB => P(4)(320),lamdaOut => P(3)(256));
U_F4257: entity F port map(lamdaA => P(4)(257),lamdaB => P(4)(321),lamdaOut => P(3)(257));
U_F4258: entity F port map(lamdaA => P(4)(258),lamdaB => P(4)(322),lamdaOut => P(3)(258));
U_F4259: entity F port map(lamdaA => P(4)(259),lamdaB => P(4)(323),lamdaOut => P(3)(259));
U_F4260: entity F port map(lamdaA => P(4)(260),lamdaB => P(4)(324),lamdaOut => P(3)(260));
U_F4261: entity F port map(lamdaA => P(4)(261),lamdaB => P(4)(325),lamdaOut => P(3)(261));
U_F4262: entity F port map(lamdaA => P(4)(262),lamdaB => P(4)(326),lamdaOut => P(3)(262));
U_F4263: entity F port map(lamdaA => P(4)(263),lamdaB => P(4)(327),lamdaOut => P(3)(263));
U_F4264: entity F port map(lamdaA => P(4)(264),lamdaB => P(4)(328),lamdaOut => P(3)(264));
U_F4265: entity F port map(lamdaA => P(4)(265),lamdaB => P(4)(329),lamdaOut => P(3)(265));
U_F4266: entity F port map(lamdaA => P(4)(266),lamdaB => P(4)(330),lamdaOut => P(3)(266));
U_F4267: entity F port map(lamdaA => P(4)(267),lamdaB => P(4)(331),lamdaOut => P(3)(267));
U_F4268: entity F port map(lamdaA => P(4)(268),lamdaB => P(4)(332),lamdaOut => P(3)(268));
U_F4269: entity F port map(lamdaA => P(4)(269),lamdaB => P(4)(333),lamdaOut => P(3)(269));
U_F4270: entity F port map(lamdaA => P(4)(270),lamdaB => P(4)(334),lamdaOut => P(3)(270));
U_F4271: entity F port map(lamdaA => P(4)(271),lamdaB => P(4)(335),lamdaOut => P(3)(271));
U_F4272: entity F port map(lamdaA => P(4)(272),lamdaB => P(4)(336),lamdaOut => P(3)(272));
U_F4273: entity F port map(lamdaA => P(4)(273),lamdaB => P(4)(337),lamdaOut => P(3)(273));
U_F4274: entity F port map(lamdaA => P(4)(274),lamdaB => P(4)(338),lamdaOut => P(3)(274));
U_F4275: entity F port map(lamdaA => P(4)(275),lamdaB => P(4)(339),lamdaOut => P(3)(275));
U_F4276: entity F port map(lamdaA => P(4)(276),lamdaB => P(4)(340),lamdaOut => P(3)(276));
U_F4277: entity F port map(lamdaA => P(4)(277),lamdaB => P(4)(341),lamdaOut => P(3)(277));
U_F4278: entity F port map(lamdaA => P(4)(278),lamdaB => P(4)(342),lamdaOut => P(3)(278));
U_F4279: entity F port map(lamdaA => P(4)(279),lamdaB => P(4)(343),lamdaOut => P(3)(279));
U_F4280: entity F port map(lamdaA => P(4)(280),lamdaB => P(4)(344),lamdaOut => P(3)(280));
U_F4281: entity F port map(lamdaA => P(4)(281),lamdaB => P(4)(345),lamdaOut => P(3)(281));
U_F4282: entity F port map(lamdaA => P(4)(282),lamdaB => P(4)(346),lamdaOut => P(3)(282));
U_F4283: entity F port map(lamdaA => P(4)(283),lamdaB => P(4)(347),lamdaOut => P(3)(283));
U_F4284: entity F port map(lamdaA => P(4)(284),lamdaB => P(4)(348),lamdaOut => P(3)(284));
U_F4285: entity F port map(lamdaA => P(4)(285),lamdaB => P(4)(349),lamdaOut => P(3)(285));
U_F4286: entity F port map(lamdaA => P(4)(286),lamdaB => P(4)(350),lamdaOut => P(3)(286));
U_F4287: entity F port map(lamdaA => P(4)(287),lamdaB => P(4)(351),lamdaOut => P(3)(287));
U_F4288: entity F port map(lamdaA => P(4)(288),lamdaB => P(4)(352),lamdaOut => P(3)(288));
U_F4289: entity F port map(lamdaA => P(4)(289),lamdaB => P(4)(353),lamdaOut => P(3)(289));
U_F4290: entity F port map(lamdaA => P(4)(290),lamdaB => P(4)(354),lamdaOut => P(3)(290));
U_F4291: entity F port map(lamdaA => P(4)(291),lamdaB => P(4)(355),lamdaOut => P(3)(291));
U_F4292: entity F port map(lamdaA => P(4)(292),lamdaB => P(4)(356),lamdaOut => P(3)(292));
U_F4293: entity F port map(lamdaA => P(4)(293),lamdaB => P(4)(357),lamdaOut => P(3)(293));
U_F4294: entity F port map(lamdaA => P(4)(294),lamdaB => P(4)(358),lamdaOut => P(3)(294));
U_F4295: entity F port map(lamdaA => P(4)(295),lamdaB => P(4)(359),lamdaOut => P(3)(295));
U_F4296: entity F port map(lamdaA => P(4)(296),lamdaB => P(4)(360),lamdaOut => P(3)(296));
U_F4297: entity F port map(lamdaA => P(4)(297),lamdaB => P(4)(361),lamdaOut => P(3)(297));
U_F4298: entity F port map(lamdaA => P(4)(298),lamdaB => P(4)(362),lamdaOut => P(3)(298));
U_F4299: entity F port map(lamdaA => P(4)(299),lamdaB => P(4)(363),lamdaOut => P(3)(299));
U_F4300: entity F port map(lamdaA => P(4)(300),lamdaB => P(4)(364),lamdaOut => P(3)(300));
U_F4301: entity F port map(lamdaA => P(4)(301),lamdaB => P(4)(365),lamdaOut => P(3)(301));
U_F4302: entity F port map(lamdaA => P(4)(302),lamdaB => P(4)(366),lamdaOut => P(3)(302));
U_F4303: entity F port map(lamdaA => P(4)(303),lamdaB => P(4)(367),lamdaOut => P(3)(303));
U_F4304: entity F port map(lamdaA => P(4)(304),lamdaB => P(4)(368),lamdaOut => P(3)(304));
U_F4305: entity F port map(lamdaA => P(4)(305),lamdaB => P(4)(369),lamdaOut => P(3)(305));
U_F4306: entity F port map(lamdaA => P(4)(306),lamdaB => P(4)(370),lamdaOut => P(3)(306));
U_F4307: entity F port map(lamdaA => P(4)(307),lamdaB => P(4)(371),lamdaOut => P(3)(307));
U_F4308: entity F port map(lamdaA => P(4)(308),lamdaB => P(4)(372),lamdaOut => P(3)(308));
U_F4309: entity F port map(lamdaA => P(4)(309),lamdaB => P(4)(373),lamdaOut => P(3)(309));
U_F4310: entity F port map(lamdaA => P(4)(310),lamdaB => P(4)(374),lamdaOut => P(3)(310));
U_F4311: entity F port map(lamdaA => P(4)(311),lamdaB => P(4)(375),lamdaOut => P(3)(311));
U_F4312: entity F port map(lamdaA => P(4)(312),lamdaB => P(4)(376),lamdaOut => P(3)(312));
U_F4313: entity F port map(lamdaA => P(4)(313),lamdaB => P(4)(377),lamdaOut => P(3)(313));
U_F4314: entity F port map(lamdaA => P(4)(314),lamdaB => P(4)(378),lamdaOut => P(3)(314));
U_F4315: entity F port map(lamdaA => P(4)(315),lamdaB => P(4)(379),lamdaOut => P(3)(315));
U_F4316: entity F port map(lamdaA => P(4)(316),lamdaB => P(4)(380),lamdaOut => P(3)(316));
U_F4317: entity F port map(lamdaA => P(4)(317),lamdaB => P(4)(381),lamdaOut => P(3)(317));
U_F4318: entity F port map(lamdaA => P(4)(318),lamdaB => P(4)(382),lamdaOut => P(3)(318));
U_F4319: entity F port map(lamdaA => P(4)(319),lamdaB => P(4)(383),lamdaOut => P(3)(319));
U_G4320: entity G port map(lamdaA => P(4)(256),lamdaB => P(4)(320),s => s(4)(128),lamdaOut => P(3)(320));
U_G4321: entity G port map(lamdaA => P(4)(257),lamdaB => P(4)(321),s => s(4)(129),lamdaOut => P(3)(321));
U_G4322: entity G port map(lamdaA => P(4)(258),lamdaB => P(4)(322),s => s(4)(130),lamdaOut => P(3)(322));
U_G4323: entity G port map(lamdaA => P(4)(259),lamdaB => P(4)(323),s => s(4)(131),lamdaOut => P(3)(323));
U_G4324: entity G port map(lamdaA => P(4)(260),lamdaB => P(4)(324),s => s(4)(132),lamdaOut => P(3)(324));
U_G4325: entity G port map(lamdaA => P(4)(261),lamdaB => P(4)(325),s => s(4)(133),lamdaOut => P(3)(325));
U_G4326: entity G port map(lamdaA => P(4)(262),lamdaB => P(4)(326),s => s(4)(134),lamdaOut => P(3)(326));
U_G4327: entity G port map(lamdaA => P(4)(263),lamdaB => P(4)(327),s => s(4)(135),lamdaOut => P(3)(327));
U_G4328: entity G port map(lamdaA => P(4)(264),lamdaB => P(4)(328),s => s(4)(136),lamdaOut => P(3)(328));
U_G4329: entity G port map(lamdaA => P(4)(265),lamdaB => P(4)(329),s => s(4)(137),lamdaOut => P(3)(329));
U_G4330: entity G port map(lamdaA => P(4)(266),lamdaB => P(4)(330),s => s(4)(138),lamdaOut => P(3)(330));
U_G4331: entity G port map(lamdaA => P(4)(267),lamdaB => P(4)(331),s => s(4)(139),lamdaOut => P(3)(331));
U_G4332: entity G port map(lamdaA => P(4)(268),lamdaB => P(4)(332),s => s(4)(140),lamdaOut => P(3)(332));
U_G4333: entity G port map(lamdaA => P(4)(269),lamdaB => P(4)(333),s => s(4)(141),lamdaOut => P(3)(333));
U_G4334: entity G port map(lamdaA => P(4)(270),lamdaB => P(4)(334),s => s(4)(142),lamdaOut => P(3)(334));
U_G4335: entity G port map(lamdaA => P(4)(271),lamdaB => P(4)(335),s => s(4)(143),lamdaOut => P(3)(335));
U_G4336: entity G port map(lamdaA => P(4)(272),lamdaB => P(4)(336),s => s(4)(144),lamdaOut => P(3)(336));
U_G4337: entity G port map(lamdaA => P(4)(273),lamdaB => P(4)(337),s => s(4)(145),lamdaOut => P(3)(337));
U_G4338: entity G port map(lamdaA => P(4)(274),lamdaB => P(4)(338),s => s(4)(146),lamdaOut => P(3)(338));
U_G4339: entity G port map(lamdaA => P(4)(275),lamdaB => P(4)(339),s => s(4)(147),lamdaOut => P(3)(339));
U_G4340: entity G port map(lamdaA => P(4)(276),lamdaB => P(4)(340),s => s(4)(148),lamdaOut => P(3)(340));
U_G4341: entity G port map(lamdaA => P(4)(277),lamdaB => P(4)(341),s => s(4)(149),lamdaOut => P(3)(341));
U_G4342: entity G port map(lamdaA => P(4)(278),lamdaB => P(4)(342),s => s(4)(150),lamdaOut => P(3)(342));
U_G4343: entity G port map(lamdaA => P(4)(279),lamdaB => P(4)(343),s => s(4)(151),lamdaOut => P(3)(343));
U_G4344: entity G port map(lamdaA => P(4)(280),lamdaB => P(4)(344),s => s(4)(152),lamdaOut => P(3)(344));
U_G4345: entity G port map(lamdaA => P(4)(281),lamdaB => P(4)(345),s => s(4)(153),lamdaOut => P(3)(345));
U_G4346: entity G port map(lamdaA => P(4)(282),lamdaB => P(4)(346),s => s(4)(154),lamdaOut => P(3)(346));
U_G4347: entity G port map(lamdaA => P(4)(283),lamdaB => P(4)(347),s => s(4)(155),lamdaOut => P(3)(347));
U_G4348: entity G port map(lamdaA => P(4)(284),lamdaB => P(4)(348),s => s(4)(156),lamdaOut => P(3)(348));
U_G4349: entity G port map(lamdaA => P(4)(285),lamdaB => P(4)(349),s => s(4)(157),lamdaOut => P(3)(349));
U_G4350: entity G port map(lamdaA => P(4)(286),lamdaB => P(4)(350),s => s(4)(158),lamdaOut => P(3)(350));
U_G4351: entity G port map(lamdaA => P(4)(287),lamdaB => P(4)(351),s => s(4)(159),lamdaOut => P(3)(351));
U_G4352: entity G port map(lamdaA => P(4)(288),lamdaB => P(4)(352),s => s(4)(160),lamdaOut => P(3)(352));
U_G4353: entity G port map(lamdaA => P(4)(289),lamdaB => P(4)(353),s => s(4)(161),lamdaOut => P(3)(353));
U_G4354: entity G port map(lamdaA => P(4)(290),lamdaB => P(4)(354),s => s(4)(162),lamdaOut => P(3)(354));
U_G4355: entity G port map(lamdaA => P(4)(291),lamdaB => P(4)(355),s => s(4)(163),lamdaOut => P(3)(355));
U_G4356: entity G port map(lamdaA => P(4)(292),lamdaB => P(4)(356),s => s(4)(164),lamdaOut => P(3)(356));
U_G4357: entity G port map(lamdaA => P(4)(293),lamdaB => P(4)(357),s => s(4)(165),lamdaOut => P(3)(357));
U_G4358: entity G port map(lamdaA => P(4)(294),lamdaB => P(4)(358),s => s(4)(166),lamdaOut => P(3)(358));
U_G4359: entity G port map(lamdaA => P(4)(295),lamdaB => P(4)(359),s => s(4)(167),lamdaOut => P(3)(359));
U_G4360: entity G port map(lamdaA => P(4)(296),lamdaB => P(4)(360),s => s(4)(168),lamdaOut => P(3)(360));
U_G4361: entity G port map(lamdaA => P(4)(297),lamdaB => P(4)(361),s => s(4)(169),lamdaOut => P(3)(361));
U_G4362: entity G port map(lamdaA => P(4)(298),lamdaB => P(4)(362),s => s(4)(170),lamdaOut => P(3)(362));
U_G4363: entity G port map(lamdaA => P(4)(299),lamdaB => P(4)(363),s => s(4)(171),lamdaOut => P(3)(363));
U_G4364: entity G port map(lamdaA => P(4)(300),lamdaB => P(4)(364),s => s(4)(172),lamdaOut => P(3)(364));
U_G4365: entity G port map(lamdaA => P(4)(301),lamdaB => P(4)(365),s => s(4)(173),lamdaOut => P(3)(365));
U_G4366: entity G port map(lamdaA => P(4)(302),lamdaB => P(4)(366),s => s(4)(174),lamdaOut => P(3)(366));
U_G4367: entity G port map(lamdaA => P(4)(303),lamdaB => P(4)(367),s => s(4)(175),lamdaOut => P(3)(367));
U_G4368: entity G port map(lamdaA => P(4)(304),lamdaB => P(4)(368),s => s(4)(176),lamdaOut => P(3)(368));
U_G4369: entity G port map(lamdaA => P(4)(305),lamdaB => P(4)(369),s => s(4)(177),lamdaOut => P(3)(369));
U_G4370: entity G port map(lamdaA => P(4)(306),lamdaB => P(4)(370),s => s(4)(178),lamdaOut => P(3)(370));
U_G4371: entity G port map(lamdaA => P(4)(307),lamdaB => P(4)(371),s => s(4)(179),lamdaOut => P(3)(371));
U_G4372: entity G port map(lamdaA => P(4)(308),lamdaB => P(4)(372),s => s(4)(180),lamdaOut => P(3)(372));
U_G4373: entity G port map(lamdaA => P(4)(309),lamdaB => P(4)(373),s => s(4)(181),lamdaOut => P(3)(373));
U_G4374: entity G port map(lamdaA => P(4)(310),lamdaB => P(4)(374),s => s(4)(182),lamdaOut => P(3)(374));
U_G4375: entity G port map(lamdaA => P(4)(311),lamdaB => P(4)(375),s => s(4)(183),lamdaOut => P(3)(375));
U_G4376: entity G port map(lamdaA => P(4)(312),lamdaB => P(4)(376),s => s(4)(184),lamdaOut => P(3)(376));
U_G4377: entity G port map(lamdaA => P(4)(313),lamdaB => P(4)(377),s => s(4)(185),lamdaOut => P(3)(377));
U_G4378: entity G port map(lamdaA => P(4)(314),lamdaB => P(4)(378),s => s(4)(186),lamdaOut => P(3)(378));
U_G4379: entity G port map(lamdaA => P(4)(315),lamdaB => P(4)(379),s => s(4)(187),lamdaOut => P(3)(379));
U_G4380: entity G port map(lamdaA => P(4)(316),lamdaB => P(4)(380),s => s(4)(188),lamdaOut => P(3)(380));
U_G4381: entity G port map(lamdaA => P(4)(317),lamdaB => P(4)(381),s => s(4)(189),lamdaOut => P(3)(381));
U_G4382: entity G port map(lamdaA => P(4)(318),lamdaB => P(4)(382),s => s(4)(190),lamdaOut => P(3)(382));
U_G4383: entity G port map(lamdaA => P(4)(319),lamdaB => P(4)(383),s => s(4)(191),lamdaOut => P(3)(383));
U_F4384: entity F port map(lamdaA => P(4)(384),lamdaB => P(4)(448),lamdaOut => P(3)(384));
U_F4385: entity F port map(lamdaA => P(4)(385),lamdaB => P(4)(449),lamdaOut => P(3)(385));
U_F4386: entity F port map(lamdaA => P(4)(386),lamdaB => P(4)(450),lamdaOut => P(3)(386));
U_F4387: entity F port map(lamdaA => P(4)(387),lamdaB => P(4)(451),lamdaOut => P(3)(387));
U_F4388: entity F port map(lamdaA => P(4)(388),lamdaB => P(4)(452),lamdaOut => P(3)(388));
U_F4389: entity F port map(lamdaA => P(4)(389),lamdaB => P(4)(453),lamdaOut => P(3)(389));
U_F4390: entity F port map(lamdaA => P(4)(390),lamdaB => P(4)(454),lamdaOut => P(3)(390));
U_F4391: entity F port map(lamdaA => P(4)(391),lamdaB => P(4)(455),lamdaOut => P(3)(391));
U_F4392: entity F port map(lamdaA => P(4)(392),lamdaB => P(4)(456),lamdaOut => P(3)(392));
U_F4393: entity F port map(lamdaA => P(4)(393),lamdaB => P(4)(457),lamdaOut => P(3)(393));
U_F4394: entity F port map(lamdaA => P(4)(394),lamdaB => P(4)(458),lamdaOut => P(3)(394));
U_F4395: entity F port map(lamdaA => P(4)(395),lamdaB => P(4)(459),lamdaOut => P(3)(395));
U_F4396: entity F port map(lamdaA => P(4)(396),lamdaB => P(4)(460),lamdaOut => P(3)(396));
U_F4397: entity F port map(lamdaA => P(4)(397),lamdaB => P(4)(461),lamdaOut => P(3)(397));
U_F4398: entity F port map(lamdaA => P(4)(398),lamdaB => P(4)(462),lamdaOut => P(3)(398));
U_F4399: entity F port map(lamdaA => P(4)(399),lamdaB => P(4)(463),lamdaOut => P(3)(399));
U_F4400: entity F port map(lamdaA => P(4)(400),lamdaB => P(4)(464),lamdaOut => P(3)(400));
U_F4401: entity F port map(lamdaA => P(4)(401),lamdaB => P(4)(465),lamdaOut => P(3)(401));
U_F4402: entity F port map(lamdaA => P(4)(402),lamdaB => P(4)(466),lamdaOut => P(3)(402));
U_F4403: entity F port map(lamdaA => P(4)(403),lamdaB => P(4)(467),lamdaOut => P(3)(403));
U_F4404: entity F port map(lamdaA => P(4)(404),lamdaB => P(4)(468),lamdaOut => P(3)(404));
U_F4405: entity F port map(lamdaA => P(4)(405),lamdaB => P(4)(469),lamdaOut => P(3)(405));
U_F4406: entity F port map(lamdaA => P(4)(406),lamdaB => P(4)(470),lamdaOut => P(3)(406));
U_F4407: entity F port map(lamdaA => P(4)(407),lamdaB => P(4)(471),lamdaOut => P(3)(407));
U_F4408: entity F port map(lamdaA => P(4)(408),lamdaB => P(4)(472),lamdaOut => P(3)(408));
U_F4409: entity F port map(lamdaA => P(4)(409),lamdaB => P(4)(473),lamdaOut => P(3)(409));
U_F4410: entity F port map(lamdaA => P(4)(410),lamdaB => P(4)(474),lamdaOut => P(3)(410));
U_F4411: entity F port map(lamdaA => P(4)(411),lamdaB => P(4)(475),lamdaOut => P(3)(411));
U_F4412: entity F port map(lamdaA => P(4)(412),lamdaB => P(4)(476),lamdaOut => P(3)(412));
U_F4413: entity F port map(lamdaA => P(4)(413),lamdaB => P(4)(477),lamdaOut => P(3)(413));
U_F4414: entity F port map(lamdaA => P(4)(414),lamdaB => P(4)(478),lamdaOut => P(3)(414));
U_F4415: entity F port map(lamdaA => P(4)(415),lamdaB => P(4)(479),lamdaOut => P(3)(415));
U_F4416: entity F port map(lamdaA => P(4)(416),lamdaB => P(4)(480),lamdaOut => P(3)(416));
U_F4417: entity F port map(lamdaA => P(4)(417),lamdaB => P(4)(481),lamdaOut => P(3)(417));
U_F4418: entity F port map(lamdaA => P(4)(418),lamdaB => P(4)(482),lamdaOut => P(3)(418));
U_F4419: entity F port map(lamdaA => P(4)(419),lamdaB => P(4)(483),lamdaOut => P(3)(419));
U_F4420: entity F port map(lamdaA => P(4)(420),lamdaB => P(4)(484),lamdaOut => P(3)(420));
U_F4421: entity F port map(lamdaA => P(4)(421),lamdaB => P(4)(485),lamdaOut => P(3)(421));
U_F4422: entity F port map(lamdaA => P(4)(422),lamdaB => P(4)(486),lamdaOut => P(3)(422));
U_F4423: entity F port map(lamdaA => P(4)(423),lamdaB => P(4)(487),lamdaOut => P(3)(423));
U_F4424: entity F port map(lamdaA => P(4)(424),lamdaB => P(4)(488),lamdaOut => P(3)(424));
U_F4425: entity F port map(lamdaA => P(4)(425),lamdaB => P(4)(489),lamdaOut => P(3)(425));
U_F4426: entity F port map(lamdaA => P(4)(426),lamdaB => P(4)(490),lamdaOut => P(3)(426));
U_F4427: entity F port map(lamdaA => P(4)(427),lamdaB => P(4)(491),lamdaOut => P(3)(427));
U_F4428: entity F port map(lamdaA => P(4)(428),lamdaB => P(4)(492),lamdaOut => P(3)(428));
U_F4429: entity F port map(lamdaA => P(4)(429),lamdaB => P(4)(493),lamdaOut => P(3)(429));
U_F4430: entity F port map(lamdaA => P(4)(430),lamdaB => P(4)(494),lamdaOut => P(3)(430));
U_F4431: entity F port map(lamdaA => P(4)(431),lamdaB => P(4)(495),lamdaOut => P(3)(431));
U_F4432: entity F port map(lamdaA => P(4)(432),lamdaB => P(4)(496),lamdaOut => P(3)(432));
U_F4433: entity F port map(lamdaA => P(4)(433),lamdaB => P(4)(497),lamdaOut => P(3)(433));
U_F4434: entity F port map(lamdaA => P(4)(434),lamdaB => P(4)(498),lamdaOut => P(3)(434));
U_F4435: entity F port map(lamdaA => P(4)(435),lamdaB => P(4)(499),lamdaOut => P(3)(435));
U_F4436: entity F port map(lamdaA => P(4)(436),lamdaB => P(4)(500),lamdaOut => P(3)(436));
U_F4437: entity F port map(lamdaA => P(4)(437),lamdaB => P(4)(501),lamdaOut => P(3)(437));
U_F4438: entity F port map(lamdaA => P(4)(438),lamdaB => P(4)(502),lamdaOut => P(3)(438));
U_F4439: entity F port map(lamdaA => P(4)(439),lamdaB => P(4)(503),lamdaOut => P(3)(439));
U_F4440: entity F port map(lamdaA => P(4)(440),lamdaB => P(4)(504),lamdaOut => P(3)(440));
U_F4441: entity F port map(lamdaA => P(4)(441),lamdaB => P(4)(505),lamdaOut => P(3)(441));
U_F4442: entity F port map(lamdaA => P(4)(442),lamdaB => P(4)(506),lamdaOut => P(3)(442));
U_F4443: entity F port map(lamdaA => P(4)(443),lamdaB => P(4)(507),lamdaOut => P(3)(443));
U_F4444: entity F port map(lamdaA => P(4)(444),lamdaB => P(4)(508),lamdaOut => P(3)(444));
U_F4445: entity F port map(lamdaA => P(4)(445),lamdaB => P(4)(509),lamdaOut => P(3)(445));
U_F4446: entity F port map(lamdaA => P(4)(446),lamdaB => P(4)(510),lamdaOut => P(3)(446));
U_F4447: entity F port map(lamdaA => P(4)(447),lamdaB => P(4)(511),lamdaOut => P(3)(447));
U_G4448: entity G port map(lamdaA => P(4)(384),lamdaB => P(4)(448),s => s(4)(192),lamdaOut => P(3)(448));
U_G4449: entity G port map(lamdaA => P(4)(385),lamdaB => P(4)(449),s => s(4)(193),lamdaOut => P(3)(449));
U_G4450: entity G port map(lamdaA => P(4)(386),lamdaB => P(4)(450),s => s(4)(194),lamdaOut => P(3)(450));
U_G4451: entity G port map(lamdaA => P(4)(387),lamdaB => P(4)(451),s => s(4)(195),lamdaOut => P(3)(451));
U_G4452: entity G port map(lamdaA => P(4)(388),lamdaB => P(4)(452),s => s(4)(196),lamdaOut => P(3)(452));
U_G4453: entity G port map(lamdaA => P(4)(389),lamdaB => P(4)(453),s => s(4)(197),lamdaOut => P(3)(453));
U_G4454: entity G port map(lamdaA => P(4)(390),lamdaB => P(4)(454),s => s(4)(198),lamdaOut => P(3)(454));
U_G4455: entity G port map(lamdaA => P(4)(391),lamdaB => P(4)(455),s => s(4)(199),lamdaOut => P(3)(455));
U_G4456: entity G port map(lamdaA => P(4)(392),lamdaB => P(4)(456),s => s(4)(200),lamdaOut => P(3)(456));
U_G4457: entity G port map(lamdaA => P(4)(393),lamdaB => P(4)(457),s => s(4)(201),lamdaOut => P(3)(457));
U_G4458: entity G port map(lamdaA => P(4)(394),lamdaB => P(4)(458),s => s(4)(202),lamdaOut => P(3)(458));
U_G4459: entity G port map(lamdaA => P(4)(395),lamdaB => P(4)(459),s => s(4)(203),lamdaOut => P(3)(459));
U_G4460: entity G port map(lamdaA => P(4)(396),lamdaB => P(4)(460),s => s(4)(204),lamdaOut => P(3)(460));
U_G4461: entity G port map(lamdaA => P(4)(397),lamdaB => P(4)(461),s => s(4)(205),lamdaOut => P(3)(461));
U_G4462: entity G port map(lamdaA => P(4)(398),lamdaB => P(4)(462),s => s(4)(206),lamdaOut => P(3)(462));
U_G4463: entity G port map(lamdaA => P(4)(399),lamdaB => P(4)(463),s => s(4)(207),lamdaOut => P(3)(463));
U_G4464: entity G port map(lamdaA => P(4)(400),lamdaB => P(4)(464),s => s(4)(208),lamdaOut => P(3)(464));
U_G4465: entity G port map(lamdaA => P(4)(401),lamdaB => P(4)(465),s => s(4)(209),lamdaOut => P(3)(465));
U_G4466: entity G port map(lamdaA => P(4)(402),lamdaB => P(4)(466),s => s(4)(210),lamdaOut => P(3)(466));
U_G4467: entity G port map(lamdaA => P(4)(403),lamdaB => P(4)(467),s => s(4)(211),lamdaOut => P(3)(467));
U_G4468: entity G port map(lamdaA => P(4)(404),lamdaB => P(4)(468),s => s(4)(212),lamdaOut => P(3)(468));
U_G4469: entity G port map(lamdaA => P(4)(405),lamdaB => P(4)(469),s => s(4)(213),lamdaOut => P(3)(469));
U_G4470: entity G port map(lamdaA => P(4)(406),lamdaB => P(4)(470),s => s(4)(214),lamdaOut => P(3)(470));
U_G4471: entity G port map(lamdaA => P(4)(407),lamdaB => P(4)(471),s => s(4)(215),lamdaOut => P(3)(471));
U_G4472: entity G port map(lamdaA => P(4)(408),lamdaB => P(4)(472),s => s(4)(216),lamdaOut => P(3)(472));
U_G4473: entity G port map(lamdaA => P(4)(409),lamdaB => P(4)(473),s => s(4)(217),lamdaOut => P(3)(473));
U_G4474: entity G port map(lamdaA => P(4)(410),lamdaB => P(4)(474),s => s(4)(218),lamdaOut => P(3)(474));
U_G4475: entity G port map(lamdaA => P(4)(411),lamdaB => P(4)(475),s => s(4)(219),lamdaOut => P(3)(475));
U_G4476: entity G port map(lamdaA => P(4)(412),lamdaB => P(4)(476),s => s(4)(220),lamdaOut => P(3)(476));
U_G4477: entity G port map(lamdaA => P(4)(413),lamdaB => P(4)(477),s => s(4)(221),lamdaOut => P(3)(477));
U_G4478: entity G port map(lamdaA => P(4)(414),lamdaB => P(4)(478),s => s(4)(222),lamdaOut => P(3)(478));
U_G4479: entity G port map(lamdaA => P(4)(415),lamdaB => P(4)(479),s => s(4)(223),lamdaOut => P(3)(479));
U_G4480: entity G port map(lamdaA => P(4)(416),lamdaB => P(4)(480),s => s(4)(224),lamdaOut => P(3)(480));
U_G4481: entity G port map(lamdaA => P(4)(417),lamdaB => P(4)(481),s => s(4)(225),lamdaOut => P(3)(481));
U_G4482: entity G port map(lamdaA => P(4)(418),lamdaB => P(4)(482),s => s(4)(226),lamdaOut => P(3)(482));
U_G4483: entity G port map(lamdaA => P(4)(419),lamdaB => P(4)(483),s => s(4)(227),lamdaOut => P(3)(483));
U_G4484: entity G port map(lamdaA => P(4)(420),lamdaB => P(4)(484),s => s(4)(228),lamdaOut => P(3)(484));
U_G4485: entity G port map(lamdaA => P(4)(421),lamdaB => P(4)(485),s => s(4)(229),lamdaOut => P(3)(485));
U_G4486: entity G port map(lamdaA => P(4)(422),lamdaB => P(4)(486),s => s(4)(230),lamdaOut => P(3)(486));
U_G4487: entity G port map(lamdaA => P(4)(423),lamdaB => P(4)(487),s => s(4)(231),lamdaOut => P(3)(487));
U_G4488: entity G port map(lamdaA => P(4)(424),lamdaB => P(4)(488),s => s(4)(232),lamdaOut => P(3)(488));
U_G4489: entity G port map(lamdaA => P(4)(425),lamdaB => P(4)(489),s => s(4)(233),lamdaOut => P(3)(489));
U_G4490: entity G port map(lamdaA => P(4)(426),lamdaB => P(4)(490),s => s(4)(234),lamdaOut => P(3)(490));
U_G4491: entity G port map(lamdaA => P(4)(427),lamdaB => P(4)(491),s => s(4)(235),lamdaOut => P(3)(491));
U_G4492: entity G port map(lamdaA => P(4)(428),lamdaB => P(4)(492),s => s(4)(236),lamdaOut => P(3)(492));
U_G4493: entity G port map(lamdaA => P(4)(429),lamdaB => P(4)(493),s => s(4)(237),lamdaOut => P(3)(493));
U_G4494: entity G port map(lamdaA => P(4)(430),lamdaB => P(4)(494),s => s(4)(238),lamdaOut => P(3)(494));
U_G4495: entity G port map(lamdaA => P(4)(431),lamdaB => P(4)(495),s => s(4)(239),lamdaOut => P(3)(495));
U_G4496: entity G port map(lamdaA => P(4)(432),lamdaB => P(4)(496),s => s(4)(240),lamdaOut => P(3)(496));
U_G4497: entity G port map(lamdaA => P(4)(433),lamdaB => P(4)(497),s => s(4)(241),lamdaOut => P(3)(497));
U_G4498: entity G port map(lamdaA => P(4)(434),lamdaB => P(4)(498),s => s(4)(242),lamdaOut => P(3)(498));
U_G4499: entity G port map(lamdaA => P(4)(435),lamdaB => P(4)(499),s => s(4)(243),lamdaOut => P(3)(499));
U_G4500: entity G port map(lamdaA => P(4)(436),lamdaB => P(4)(500),s => s(4)(244),lamdaOut => P(3)(500));
U_G4501: entity G port map(lamdaA => P(4)(437),lamdaB => P(4)(501),s => s(4)(245),lamdaOut => P(3)(501));
U_G4502: entity G port map(lamdaA => P(4)(438),lamdaB => P(4)(502),s => s(4)(246),lamdaOut => P(3)(502));
U_G4503: entity G port map(lamdaA => P(4)(439),lamdaB => P(4)(503),s => s(4)(247),lamdaOut => P(3)(503));
U_G4504: entity G port map(lamdaA => P(4)(440),lamdaB => P(4)(504),s => s(4)(248),lamdaOut => P(3)(504));
U_G4505: entity G port map(lamdaA => P(4)(441),lamdaB => P(4)(505),s => s(4)(249),lamdaOut => P(3)(505));
U_G4506: entity G port map(lamdaA => P(4)(442),lamdaB => P(4)(506),s => s(4)(250),lamdaOut => P(3)(506));
U_G4507: entity G port map(lamdaA => P(4)(443),lamdaB => P(4)(507),s => s(4)(251),lamdaOut => P(3)(507));
U_G4508: entity G port map(lamdaA => P(4)(444),lamdaB => P(4)(508),s => s(4)(252),lamdaOut => P(3)(508));
U_G4509: entity G port map(lamdaA => P(4)(445),lamdaB => P(4)(509),s => s(4)(253),lamdaOut => P(3)(509));
U_G4510: entity G port map(lamdaA => P(4)(446),lamdaB => P(4)(510),s => s(4)(254),lamdaOut => P(3)(510));
U_G4511: entity G port map(lamdaA => P(4)(447),lamdaB => P(4)(511),s => s(4)(255),lamdaOut => P(3)(511));
U_F4512: entity F port map(lamdaA => P(4)(512),lamdaB => P(4)(576),lamdaOut => P(3)(512));
U_F4513: entity F port map(lamdaA => P(4)(513),lamdaB => P(4)(577),lamdaOut => P(3)(513));
U_F4514: entity F port map(lamdaA => P(4)(514),lamdaB => P(4)(578),lamdaOut => P(3)(514));
U_F4515: entity F port map(lamdaA => P(4)(515),lamdaB => P(4)(579),lamdaOut => P(3)(515));
U_F4516: entity F port map(lamdaA => P(4)(516),lamdaB => P(4)(580),lamdaOut => P(3)(516));
U_F4517: entity F port map(lamdaA => P(4)(517),lamdaB => P(4)(581),lamdaOut => P(3)(517));
U_F4518: entity F port map(lamdaA => P(4)(518),lamdaB => P(4)(582),lamdaOut => P(3)(518));
U_F4519: entity F port map(lamdaA => P(4)(519),lamdaB => P(4)(583),lamdaOut => P(3)(519));
U_F4520: entity F port map(lamdaA => P(4)(520),lamdaB => P(4)(584),lamdaOut => P(3)(520));
U_F4521: entity F port map(lamdaA => P(4)(521),lamdaB => P(4)(585),lamdaOut => P(3)(521));
U_F4522: entity F port map(lamdaA => P(4)(522),lamdaB => P(4)(586),lamdaOut => P(3)(522));
U_F4523: entity F port map(lamdaA => P(4)(523),lamdaB => P(4)(587),lamdaOut => P(3)(523));
U_F4524: entity F port map(lamdaA => P(4)(524),lamdaB => P(4)(588),lamdaOut => P(3)(524));
U_F4525: entity F port map(lamdaA => P(4)(525),lamdaB => P(4)(589),lamdaOut => P(3)(525));
U_F4526: entity F port map(lamdaA => P(4)(526),lamdaB => P(4)(590),lamdaOut => P(3)(526));
U_F4527: entity F port map(lamdaA => P(4)(527),lamdaB => P(4)(591),lamdaOut => P(3)(527));
U_F4528: entity F port map(lamdaA => P(4)(528),lamdaB => P(4)(592),lamdaOut => P(3)(528));
U_F4529: entity F port map(lamdaA => P(4)(529),lamdaB => P(4)(593),lamdaOut => P(3)(529));
U_F4530: entity F port map(lamdaA => P(4)(530),lamdaB => P(4)(594),lamdaOut => P(3)(530));
U_F4531: entity F port map(lamdaA => P(4)(531),lamdaB => P(4)(595),lamdaOut => P(3)(531));
U_F4532: entity F port map(lamdaA => P(4)(532),lamdaB => P(4)(596),lamdaOut => P(3)(532));
U_F4533: entity F port map(lamdaA => P(4)(533),lamdaB => P(4)(597),lamdaOut => P(3)(533));
U_F4534: entity F port map(lamdaA => P(4)(534),lamdaB => P(4)(598),lamdaOut => P(3)(534));
U_F4535: entity F port map(lamdaA => P(4)(535),lamdaB => P(4)(599),lamdaOut => P(3)(535));
U_F4536: entity F port map(lamdaA => P(4)(536),lamdaB => P(4)(600),lamdaOut => P(3)(536));
U_F4537: entity F port map(lamdaA => P(4)(537),lamdaB => P(4)(601),lamdaOut => P(3)(537));
U_F4538: entity F port map(lamdaA => P(4)(538),lamdaB => P(4)(602),lamdaOut => P(3)(538));
U_F4539: entity F port map(lamdaA => P(4)(539),lamdaB => P(4)(603),lamdaOut => P(3)(539));
U_F4540: entity F port map(lamdaA => P(4)(540),lamdaB => P(4)(604),lamdaOut => P(3)(540));
U_F4541: entity F port map(lamdaA => P(4)(541),lamdaB => P(4)(605),lamdaOut => P(3)(541));
U_F4542: entity F port map(lamdaA => P(4)(542),lamdaB => P(4)(606),lamdaOut => P(3)(542));
U_F4543: entity F port map(lamdaA => P(4)(543),lamdaB => P(4)(607),lamdaOut => P(3)(543));
U_F4544: entity F port map(lamdaA => P(4)(544),lamdaB => P(4)(608),lamdaOut => P(3)(544));
U_F4545: entity F port map(lamdaA => P(4)(545),lamdaB => P(4)(609),lamdaOut => P(3)(545));
U_F4546: entity F port map(lamdaA => P(4)(546),lamdaB => P(4)(610),lamdaOut => P(3)(546));
U_F4547: entity F port map(lamdaA => P(4)(547),lamdaB => P(4)(611),lamdaOut => P(3)(547));
U_F4548: entity F port map(lamdaA => P(4)(548),lamdaB => P(4)(612),lamdaOut => P(3)(548));
U_F4549: entity F port map(lamdaA => P(4)(549),lamdaB => P(4)(613),lamdaOut => P(3)(549));
U_F4550: entity F port map(lamdaA => P(4)(550),lamdaB => P(4)(614),lamdaOut => P(3)(550));
U_F4551: entity F port map(lamdaA => P(4)(551),lamdaB => P(4)(615),lamdaOut => P(3)(551));
U_F4552: entity F port map(lamdaA => P(4)(552),lamdaB => P(4)(616),lamdaOut => P(3)(552));
U_F4553: entity F port map(lamdaA => P(4)(553),lamdaB => P(4)(617),lamdaOut => P(3)(553));
U_F4554: entity F port map(lamdaA => P(4)(554),lamdaB => P(4)(618),lamdaOut => P(3)(554));
U_F4555: entity F port map(lamdaA => P(4)(555),lamdaB => P(4)(619),lamdaOut => P(3)(555));
U_F4556: entity F port map(lamdaA => P(4)(556),lamdaB => P(4)(620),lamdaOut => P(3)(556));
U_F4557: entity F port map(lamdaA => P(4)(557),lamdaB => P(4)(621),lamdaOut => P(3)(557));
U_F4558: entity F port map(lamdaA => P(4)(558),lamdaB => P(4)(622),lamdaOut => P(3)(558));
U_F4559: entity F port map(lamdaA => P(4)(559),lamdaB => P(4)(623),lamdaOut => P(3)(559));
U_F4560: entity F port map(lamdaA => P(4)(560),lamdaB => P(4)(624),lamdaOut => P(3)(560));
U_F4561: entity F port map(lamdaA => P(4)(561),lamdaB => P(4)(625),lamdaOut => P(3)(561));
U_F4562: entity F port map(lamdaA => P(4)(562),lamdaB => P(4)(626),lamdaOut => P(3)(562));
U_F4563: entity F port map(lamdaA => P(4)(563),lamdaB => P(4)(627),lamdaOut => P(3)(563));
U_F4564: entity F port map(lamdaA => P(4)(564),lamdaB => P(4)(628),lamdaOut => P(3)(564));
U_F4565: entity F port map(lamdaA => P(4)(565),lamdaB => P(4)(629),lamdaOut => P(3)(565));
U_F4566: entity F port map(lamdaA => P(4)(566),lamdaB => P(4)(630),lamdaOut => P(3)(566));
U_F4567: entity F port map(lamdaA => P(4)(567),lamdaB => P(4)(631),lamdaOut => P(3)(567));
U_F4568: entity F port map(lamdaA => P(4)(568),lamdaB => P(4)(632),lamdaOut => P(3)(568));
U_F4569: entity F port map(lamdaA => P(4)(569),lamdaB => P(4)(633),lamdaOut => P(3)(569));
U_F4570: entity F port map(lamdaA => P(4)(570),lamdaB => P(4)(634),lamdaOut => P(3)(570));
U_F4571: entity F port map(lamdaA => P(4)(571),lamdaB => P(4)(635),lamdaOut => P(3)(571));
U_F4572: entity F port map(lamdaA => P(4)(572),lamdaB => P(4)(636),lamdaOut => P(3)(572));
U_F4573: entity F port map(lamdaA => P(4)(573),lamdaB => P(4)(637),lamdaOut => P(3)(573));
U_F4574: entity F port map(lamdaA => P(4)(574),lamdaB => P(4)(638),lamdaOut => P(3)(574));
U_F4575: entity F port map(lamdaA => P(4)(575),lamdaB => P(4)(639),lamdaOut => P(3)(575));
U_G4576: entity G port map(lamdaA => P(4)(512),lamdaB => P(4)(576),s => s(4)(256),lamdaOut => P(3)(576));
U_G4577: entity G port map(lamdaA => P(4)(513),lamdaB => P(4)(577),s => s(4)(257),lamdaOut => P(3)(577));
U_G4578: entity G port map(lamdaA => P(4)(514),lamdaB => P(4)(578),s => s(4)(258),lamdaOut => P(3)(578));
U_G4579: entity G port map(lamdaA => P(4)(515),lamdaB => P(4)(579),s => s(4)(259),lamdaOut => P(3)(579));
U_G4580: entity G port map(lamdaA => P(4)(516),lamdaB => P(4)(580),s => s(4)(260),lamdaOut => P(3)(580));
U_G4581: entity G port map(lamdaA => P(4)(517),lamdaB => P(4)(581),s => s(4)(261),lamdaOut => P(3)(581));
U_G4582: entity G port map(lamdaA => P(4)(518),lamdaB => P(4)(582),s => s(4)(262),lamdaOut => P(3)(582));
U_G4583: entity G port map(lamdaA => P(4)(519),lamdaB => P(4)(583),s => s(4)(263),lamdaOut => P(3)(583));
U_G4584: entity G port map(lamdaA => P(4)(520),lamdaB => P(4)(584),s => s(4)(264),lamdaOut => P(3)(584));
U_G4585: entity G port map(lamdaA => P(4)(521),lamdaB => P(4)(585),s => s(4)(265),lamdaOut => P(3)(585));
U_G4586: entity G port map(lamdaA => P(4)(522),lamdaB => P(4)(586),s => s(4)(266),lamdaOut => P(3)(586));
U_G4587: entity G port map(lamdaA => P(4)(523),lamdaB => P(4)(587),s => s(4)(267),lamdaOut => P(3)(587));
U_G4588: entity G port map(lamdaA => P(4)(524),lamdaB => P(4)(588),s => s(4)(268),lamdaOut => P(3)(588));
U_G4589: entity G port map(lamdaA => P(4)(525),lamdaB => P(4)(589),s => s(4)(269),lamdaOut => P(3)(589));
U_G4590: entity G port map(lamdaA => P(4)(526),lamdaB => P(4)(590),s => s(4)(270),lamdaOut => P(3)(590));
U_G4591: entity G port map(lamdaA => P(4)(527),lamdaB => P(4)(591),s => s(4)(271),lamdaOut => P(3)(591));
U_G4592: entity G port map(lamdaA => P(4)(528),lamdaB => P(4)(592),s => s(4)(272),lamdaOut => P(3)(592));
U_G4593: entity G port map(lamdaA => P(4)(529),lamdaB => P(4)(593),s => s(4)(273),lamdaOut => P(3)(593));
U_G4594: entity G port map(lamdaA => P(4)(530),lamdaB => P(4)(594),s => s(4)(274),lamdaOut => P(3)(594));
U_G4595: entity G port map(lamdaA => P(4)(531),lamdaB => P(4)(595),s => s(4)(275),lamdaOut => P(3)(595));
U_G4596: entity G port map(lamdaA => P(4)(532),lamdaB => P(4)(596),s => s(4)(276),lamdaOut => P(3)(596));
U_G4597: entity G port map(lamdaA => P(4)(533),lamdaB => P(4)(597),s => s(4)(277),lamdaOut => P(3)(597));
U_G4598: entity G port map(lamdaA => P(4)(534),lamdaB => P(4)(598),s => s(4)(278),lamdaOut => P(3)(598));
U_G4599: entity G port map(lamdaA => P(4)(535),lamdaB => P(4)(599),s => s(4)(279),lamdaOut => P(3)(599));
U_G4600: entity G port map(lamdaA => P(4)(536),lamdaB => P(4)(600),s => s(4)(280),lamdaOut => P(3)(600));
U_G4601: entity G port map(lamdaA => P(4)(537),lamdaB => P(4)(601),s => s(4)(281),lamdaOut => P(3)(601));
U_G4602: entity G port map(lamdaA => P(4)(538),lamdaB => P(4)(602),s => s(4)(282),lamdaOut => P(3)(602));
U_G4603: entity G port map(lamdaA => P(4)(539),lamdaB => P(4)(603),s => s(4)(283),lamdaOut => P(3)(603));
U_G4604: entity G port map(lamdaA => P(4)(540),lamdaB => P(4)(604),s => s(4)(284),lamdaOut => P(3)(604));
U_G4605: entity G port map(lamdaA => P(4)(541),lamdaB => P(4)(605),s => s(4)(285),lamdaOut => P(3)(605));
U_G4606: entity G port map(lamdaA => P(4)(542),lamdaB => P(4)(606),s => s(4)(286),lamdaOut => P(3)(606));
U_G4607: entity G port map(lamdaA => P(4)(543),lamdaB => P(4)(607),s => s(4)(287),lamdaOut => P(3)(607));
U_G4608: entity G port map(lamdaA => P(4)(544),lamdaB => P(4)(608),s => s(4)(288),lamdaOut => P(3)(608));
U_G4609: entity G port map(lamdaA => P(4)(545),lamdaB => P(4)(609),s => s(4)(289),lamdaOut => P(3)(609));
U_G4610: entity G port map(lamdaA => P(4)(546),lamdaB => P(4)(610),s => s(4)(290),lamdaOut => P(3)(610));
U_G4611: entity G port map(lamdaA => P(4)(547),lamdaB => P(4)(611),s => s(4)(291),lamdaOut => P(3)(611));
U_G4612: entity G port map(lamdaA => P(4)(548),lamdaB => P(4)(612),s => s(4)(292),lamdaOut => P(3)(612));
U_G4613: entity G port map(lamdaA => P(4)(549),lamdaB => P(4)(613),s => s(4)(293),lamdaOut => P(3)(613));
U_G4614: entity G port map(lamdaA => P(4)(550),lamdaB => P(4)(614),s => s(4)(294),lamdaOut => P(3)(614));
U_G4615: entity G port map(lamdaA => P(4)(551),lamdaB => P(4)(615),s => s(4)(295),lamdaOut => P(3)(615));
U_G4616: entity G port map(lamdaA => P(4)(552),lamdaB => P(4)(616),s => s(4)(296),lamdaOut => P(3)(616));
U_G4617: entity G port map(lamdaA => P(4)(553),lamdaB => P(4)(617),s => s(4)(297),lamdaOut => P(3)(617));
U_G4618: entity G port map(lamdaA => P(4)(554),lamdaB => P(4)(618),s => s(4)(298),lamdaOut => P(3)(618));
U_G4619: entity G port map(lamdaA => P(4)(555),lamdaB => P(4)(619),s => s(4)(299),lamdaOut => P(3)(619));
U_G4620: entity G port map(lamdaA => P(4)(556),lamdaB => P(4)(620),s => s(4)(300),lamdaOut => P(3)(620));
U_G4621: entity G port map(lamdaA => P(4)(557),lamdaB => P(4)(621),s => s(4)(301),lamdaOut => P(3)(621));
U_G4622: entity G port map(lamdaA => P(4)(558),lamdaB => P(4)(622),s => s(4)(302),lamdaOut => P(3)(622));
U_G4623: entity G port map(lamdaA => P(4)(559),lamdaB => P(4)(623),s => s(4)(303),lamdaOut => P(3)(623));
U_G4624: entity G port map(lamdaA => P(4)(560),lamdaB => P(4)(624),s => s(4)(304),lamdaOut => P(3)(624));
U_G4625: entity G port map(lamdaA => P(4)(561),lamdaB => P(4)(625),s => s(4)(305),lamdaOut => P(3)(625));
U_G4626: entity G port map(lamdaA => P(4)(562),lamdaB => P(4)(626),s => s(4)(306),lamdaOut => P(3)(626));
U_G4627: entity G port map(lamdaA => P(4)(563),lamdaB => P(4)(627),s => s(4)(307),lamdaOut => P(3)(627));
U_G4628: entity G port map(lamdaA => P(4)(564),lamdaB => P(4)(628),s => s(4)(308),lamdaOut => P(3)(628));
U_G4629: entity G port map(lamdaA => P(4)(565),lamdaB => P(4)(629),s => s(4)(309),lamdaOut => P(3)(629));
U_G4630: entity G port map(lamdaA => P(4)(566),lamdaB => P(4)(630),s => s(4)(310),lamdaOut => P(3)(630));
U_G4631: entity G port map(lamdaA => P(4)(567),lamdaB => P(4)(631),s => s(4)(311),lamdaOut => P(3)(631));
U_G4632: entity G port map(lamdaA => P(4)(568),lamdaB => P(4)(632),s => s(4)(312),lamdaOut => P(3)(632));
U_G4633: entity G port map(lamdaA => P(4)(569),lamdaB => P(4)(633),s => s(4)(313),lamdaOut => P(3)(633));
U_G4634: entity G port map(lamdaA => P(4)(570),lamdaB => P(4)(634),s => s(4)(314),lamdaOut => P(3)(634));
U_G4635: entity G port map(lamdaA => P(4)(571),lamdaB => P(4)(635),s => s(4)(315),lamdaOut => P(3)(635));
U_G4636: entity G port map(lamdaA => P(4)(572),lamdaB => P(4)(636),s => s(4)(316),lamdaOut => P(3)(636));
U_G4637: entity G port map(lamdaA => P(4)(573),lamdaB => P(4)(637),s => s(4)(317),lamdaOut => P(3)(637));
U_G4638: entity G port map(lamdaA => P(4)(574),lamdaB => P(4)(638),s => s(4)(318),lamdaOut => P(3)(638));
U_G4639: entity G port map(lamdaA => P(4)(575),lamdaB => P(4)(639),s => s(4)(319),lamdaOut => P(3)(639));
U_F4640: entity F port map(lamdaA => P(4)(640),lamdaB => P(4)(704),lamdaOut => P(3)(640));
U_F4641: entity F port map(lamdaA => P(4)(641),lamdaB => P(4)(705),lamdaOut => P(3)(641));
U_F4642: entity F port map(lamdaA => P(4)(642),lamdaB => P(4)(706),lamdaOut => P(3)(642));
U_F4643: entity F port map(lamdaA => P(4)(643),lamdaB => P(4)(707),lamdaOut => P(3)(643));
U_F4644: entity F port map(lamdaA => P(4)(644),lamdaB => P(4)(708),lamdaOut => P(3)(644));
U_F4645: entity F port map(lamdaA => P(4)(645),lamdaB => P(4)(709),lamdaOut => P(3)(645));
U_F4646: entity F port map(lamdaA => P(4)(646),lamdaB => P(4)(710),lamdaOut => P(3)(646));
U_F4647: entity F port map(lamdaA => P(4)(647),lamdaB => P(4)(711),lamdaOut => P(3)(647));
U_F4648: entity F port map(lamdaA => P(4)(648),lamdaB => P(4)(712),lamdaOut => P(3)(648));
U_F4649: entity F port map(lamdaA => P(4)(649),lamdaB => P(4)(713),lamdaOut => P(3)(649));
U_F4650: entity F port map(lamdaA => P(4)(650),lamdaB => P(4)(714),lamdaOut => P(3)(650));
U_F4651: entity F port map(lamdaA => P(4)(651),lamdaB => P(4)(715),lamdaOut => P(3)(651));
U_F4652: entity F port map(lamdaA => P(4)(652),lamdaB => P(4)(716),lamdaOut => P(3)(652));
U_F4653: entity F port map(lamdaA => P(4)(653),lamdaB => P(4)(717),lamdaOut => P(3)(653));
U_F4654: entity F port map(lamdaA => P(4)(654),lamdaB => P(4)(718),lamdaOut => P(3)(654));
U_F4655: entity F port map(lamdaA => P(4)(655),lamdaB => P(4)(719),lamdaOut => P(3)(655));
U_F4656: entity F port map(lamdaA => P(4)(656),lamdaB => P(4)(720),lamdaOut => P(3)(656));
U_F4657: entity F port map(lamdaA => P(4)(657),lamdaB => P(4)(721),lamdaOut => P(3)(657));
U_F4658: entity F port map(lamdaA => P(4)(658),lamdaB => P(4)(722),lamdaOut => P(3)(658));
U_F4659: entity F port map(lamdaA => P(4)(659),lamdaB => P(4)(723),lamdaOut => P(3)(659));
U_F4660: entity F port map(lamdaA => P(4)(660),lamdaB => P(4)(724),lamdaOut => P(3)(660));
U_F4661: entity F port map(lamdaA => P(4)(661),lamdaB => P(4)(725),lamdaOut => P(3)(661));
U_F4662: entity F port map(lamdaA => P(4)(662),lamdaB => P(4)(726),lamdaOut => P(3)(662));
U_F4663: entity F port map(lamdaA => P(4)(663),lamdaB => P(4)(727),lamdaOut => P(3)(663));
U_F4664: entity F port map(lamdaA => P(4)(664),lamdaB => P(4)(728),lamdaOut => P(3)(664));
U_F4665: entity F port map(lamdaA => P(4)(665),lamdaB => P(4)(729),lamdaOut => P(3)(665));
U_F4666: entity F port map(lamdaA => P(4)(666),lamdaB => P(4)(730),lamdaOut => P(3)(666));
U_F4667: entity F port map(lamdaA => P(4)(667),lamdaB => P(4)(731),lamdaOut => P(3)(667));
U_F4668: entity F port map(lamdaA => P(4)(668),lamdaB => P(4)(732),lamdaOut => P(3)(668));
U_F4669: entity F port map(lamdaA => P(4)(669),lamdaB => P(4)(733),lamdaOut => P(3)(669));
U_F4670: entity F port map(lamdaA => P(4)(670),lamdaB => P(4)(734),lamdaOut => P(3)(670));
U_F4671: entity F port map(lamdaA => P(4)(671),lamdaB => P(4)(735),lamdaOut => P(3)(671));
U_F4672: entity F port map(lamdaA => P(4)(672),lamdaB => P(4)(736),lamdaOut => P(3)(672));
U_F4673: entity F port map(lamdaA => P(4)(673),lamdaB => P(4)(737),lamdaOut => P(3)(673));
U_F4674: entity F port map(lamdaA => P(4)(674),lamdaB => P(4)(738),lamdaOut => P(3)(674));
U_F4675: entity F port map(lamdaA => P(4)(675),lamdaB => P(4)(739),lamdaOut => P(3)(675));
U_F4676: entity F port map(lamdaA => P(4)(676),lamdaB => P(4)(740),lamdaOut => P(3)(676));
U_F4677: entity F port map(lamdaA => P(4)(677),lamdaB => P(4)(741),lamdaOut => P(3)(677));
U_F4678: entity F port map(lamdaA => P(4)(678),lamdaB => P(4)(742),lamdaOut => P(3)(678));
U_F4679: entity F port map(lamdaA => P(4)(679),lamdaB => P(4)(743),lamdaOut => P(3)(679));
U_F4680: entity F port map(lamdaA => P(4)(680),lamdaB => P(4)(744),lamdaOut => P(3)(680));
U_F4681: entity F port map(lamdaA => P(4)(681),lamdaB => P(4)(745),lamdaOut => P(3)(681));
U_F4682: entity F port map(lamdaA => P(4)(682),lamdaB => P(4)(746),lamdaOut => P(3)(682));
U_F4683: entity F port map(lamdaA => P(4)(683),lamdaB => P(4)(747),lamdaOut => P(3)(683));
U_F4684: entity F port map(lamdaA => P(4)(684),lamdaB => P(4)(748),lamdaOut => P(3)(684));
U_F4685: entity F port map(lamdaA => P(4)(685),lamdaB => P(4)(749),lamdaOut => P(3)(685));
U_F4686: entity F port map(lamdaA => P(4)(686),lamdaB => P(4)(750),lamdaOut => P(3)(686));
U_F4687: entity F port map(lamdaA => P(4)(687),lamdaB => P(4)(751),lamdaOut => P(3)(687));
U_F4688: entity F port map(lamdaA => P(4)(688),lamdaB => P(4)(752),lamdaOut => P(3)(688));
U_F4689: entity F port map(lamdaA => P(4)(689),lamdaB => P(4)(753),lamdaOut => P(3)(689));
U_F4690: entity F port map(lamdaA => P(4)(690),lamdaB => P(4)(754),lamdaOut => P(3)(690));
U_F4691: entity F port map(lamdaA => P(4)(691),lamdaB => P(4)(755),lamdaOut => P(3)(691));
U_F4692: entity F port map(lamdaA => P(4)(692),lamdaB => P(4)(756),lamdaOut => P(3)(692));
U_F4693: entity F port map(lamdaA => P(4)(693),lamdaB => P(4)(757),lamdaOut => P(3)(693));
U_F4694: entity F port map(lamdaA => P(4)(694),lamdaB => P(4)(758),lamdaOut => P(3)(694));
U_F4695: entity F port map(lamdaA => P(4)(695),lamdaB => P(4)(759),lamdaOut => P(3)(695));
U_F4696: entity F port map(lamdaA => P(4)(696),lamdaB => P(4)(760),lamdaOut => P(3)(696));
U_F4697: entity F port map(lamdaA => P(4)(697),lamdaB => P(4)(761),lamdaOut => P(3)(697));
U_F4698: entity F port map(lamdaA => P(4)(698),lamdaB => P(4)(762),lamdaOut => P(3)(698));
U_F4699: entity F port map(lamdaA => P(4)(699),lamdaB => P(4)(763),lamdaOut => P(3)(699));
U_F4700: entity F port map(lamdaA => P(4)(700),lamdaB => P(4)(764),lamdaOut => P(3)(700));
U_F4701: entity F port map(lamdaA => P(4)(701),lamdaB => P(4)(765),lamdaOut => P(3)(701));
U_F4702: entity F port map(lamdaA => P(4)(702),lamdaB => P(4)(766),lamdaOut => P(3)(702));
U_F4703: entity F port map(lamdaA => P(4)(703),lamdaB => P(4)(767),lamdaOut => P(3)(703));
U_G4704: entity G port map(lamdaA => P(4)(640),lamdaB => P(4)(704),s => s(4)(320),lamdaOut => P(3)(704));
U_G4705: entity G port map(lamdaA => P(4)(641),lamdaB => P(4)(705),s => s(4)(321),lamdaOut => P(3)(705));
U_G4706: entity G port map(lamdaA => P(4)(642),lamdaB => P(4)(706),s => s(4)(322),lamdaOut => P(3)(706));
U_G4707: entity G port map(lamdaA => P(4)(643),lamdaB => P(4)(707),s => s(4)(323),lamdaOut => P(3)(707));
U_G4708: entity G port map(lamdaA => P(4)(644),lamdaB => P(4)(708),s => s(4)(324),lamdaOut => P(3)(708));
U_G4709: entity G port map(lamdaA => P(4)(645),lamdaB => P(4)(709),s => s(4)(325),lamdaOut => P(3)(709));
U_G4710: entity G port map(lamdaA => P(4)(646),lamdaB => P(4)(710),s => s(4)(326),lamdaOut => P(3)(710));
U_G4711: entity G port map(lamdaA => P(4)(647),lamdaB => P(4)(711),s => s(4)(327),lamdaOut => P(3)(711));
U_G4712: entity G port map(lamdaA => P(4)(648),lamdaB => P(4)(712),s => s(4)(328),lamdaOut => P(3)(712));
U_G4713: entity G port map(lamdaA => P(4)(649),lamdaB => P(4)(713),s => s(4)(329),lamdaOut => P(3)(713));
U_G4714: entity G port map(lamdaA => P(4)(650),lamdaB => P(4)(714),s => s(4)(330),lamdaOut => P(3)(714));
U_G4715: entity G port map(lamdaA => P(4)(651),lamdaB => P(4)(715),s => s(4)(331),lamdaOut => P(3)(715));
U_G4716: entity G port map(lamdaA => P(4)(652),lamdaB => P(4)(716),s => s(4)(332),lamdaOut => P(3)(716));
U_G4717: entity G port map(lamdaA => P(4)(653),lamdaB => P(4)(717),s => s(4)(333),lamdaOut => P(3)(717));
U_G4718: entity G port map(lamdaA => P(4)(654),lamdaB => P(4)(718),s => s(4)(334),lamdaOut => P(3)(718));
U_G4719: entity G port map(lamdaA => P(4)(655),lamdaB => P(4)(719),s => s(4)(335),lamdaOut => P(3)(719));
U_G4720: entity G port map(lamdaA => P(4)(656),lamdaB => P(4)(720),s => s(4)(336),lamdaOut => P(3)(720));
U_G4721: entity G port map(lamdaA => P(4)(657),lamdaB => P(4)(721),s => s(4)(337),lamdaOut => P(3)(721));
U_G4722: entity G port map(lamdaA => P(4)(658),lamdaB => P(4)(722),s => s(4)(338),lamdaOut => P(3)(722));
U_G4723: entity G port map(lamdaA => P(4)(659),lamdaB => P(4)(723),s => s(4)(339),lamdaOut => P(3)(723));
U_G4724: entity G port map(lamdaA => P(4)(660),lamdaB => P(4)(724),s => s(4)(340),lamdaOut => P(3)(724));
U_G4725: entity G port map(lamdaA => P(4)(661),lamdaB => P(4)(725),s => s(4)(341),lamdaOut => P(3)(725));
U_G4726: entity G port map(lamdaA => P(4)(662),lamdaB => P(4)(726),s => s(4)(342),lamdaOut => P(3)(726));
U_G4727: entity G port map(lamdaA => P(4)(663),lamdaB => P(4)(727),s => s(4)(343),lamdaOut => P(3)(727));
U_G4728: entity G port map(lamdaA => P(4)(664),lamdaB => P(4)(728),s => s(4)(344),lamdaOut => P(3)(728));
U_G4729: entity G port map(lamdaA => P(4)(665),lamdaB => P(4)(729),s => s(4)(345),lamdaOut => P(3)(729));
U_G4730: entity G port map(lamdaA => P(4)(666),lamdaB => P(4)(730),s => s(4)(346),lamdaOut => P(3)(730));
U_G4731: entity G port map(lamdaA => P(4)(667),lamdaB => P(4)(731),s => s(4)(347),lamdaOut => P(3)(731));
U_G4732: entity G port map(lamdaA => P(4)(668),lamdaB => P(4)(732),s => s(4)(348),lamdaOut => P(3)(732));
U_G4733: entity G port map(lamdaA => P(4)(669),lamdaB => P(4)(733),s => s(4)(349),lamdaOut => P(3)(733));
U_G4734: entity G port map(lamdaA => P(4)(670),lamdaB => P(4)(734),s => s(4)(350),lamdaOut => P(3)(734));
U_G4735: entity G port map(lamdaA => P(4)(671),lamdaB => P(4)(735),s => s(4)(351),lamdaOut => P(3)(735));
U_G4736: entity G port map(lamdaA => P(4)(672),lamdaB => P(4)(736),s => s(4)(352),lamdaOut => P(3)(736));
U_G4737: entity G port map(lamdaA => P(4)(673),lamdaB => P(4)(737),s => s(4)(353),lamdaOut => P(3)(737));
U_G4738: entity G port map(lamdaA => P(4)(674),lamdaB => P(4)(738),s => s(4)(354),lamdaOut => P(3)(738));
U_G4739: entity G port map(lamdaA => P(4)(675),lamdaB => P(4)(739),s => s(4)(355),lamdaOut => P(3)(739));
U_G4740: entity G port map(lamdaA => P(4)(676),lamdaB => P(4)(740),s => s(4)(356),lamdaOut => P(3)(740));
U_G4741: entity G port map(lamdaA => P(4)(677),lamdaB => P(4)(741),s => s(4)(357),lamdaOut => P(3)(741));
U_G4742: entity G port map(lamdaA => P(4)(678),lamdaB => P(4)(742),s => s(4)(358),lamdaOut => P(3)(742));
U_G4743: entity G port map(lamdaA => P(4)(679),lamdaB => P(4)(743),s => s(4)(359),lamdaOut => P(3)(743));
U_G4744: entity G port map(lamdaA => P(4)(680),lamdaB => P(4)(744),s => s(4)(360),lamdaOut => P(3)(744));
U_G4745: entity G port map(lamdaA => P(4)(681),lamdaB => P(4)(745),s => s(4)(361),lamdaOut => P(3)(745));
U_G4746: entity G port map(lamdaA => P(4)(682),lamdaB => P(4)(746),s => s(4)(362),lamdaOut => P(3)(746));
U_G4747: entity G port map(lamdaA => P(4)(683),lamdaB => P(4)(747),s => s(4)(363),lamdaOut => P(3)(747));
U_G4748: entity G port map(lamdaA => P(4)(684),lamdaB => P(4)(748),s => s(4)(364),lamdaOut => P(3)(748));
U_G4749: entity G port map(lamdaA => P(4)(685),lamdaB => P(4)(749),s => s(4)(365),lamdaOut => P(3)(749));
U_G4750: entity G port map(lamdaA => P(4)(686),lamdaB => P(4)(750),s => s(4)(366),lamdaOut => P(3)(750));
U_G4751: entity G port map(lamdaA => P(4)(687),lamdaB => P(4)(751),s => s(4)(367),lamdaOut => P(3)(751));
U_G4752: entity G port map(lamdaA => P(4)(688),lamdaB => P(4)(752),s => s(4)(368),lamdaOut => P(3)(752));
U_G4753: entity G port map(lamdaA => P(4)(689),lamdaB => P(4)(753),s => s(4)(369),lamdaOut => P(3)(753));
U_G4754: entity G port map(lamdaA => P(4)(690),lamdaB => P(4)(754),s => s(4)(370),lamdaOut => P(3)(754));
U_G4755: entity G port map(lamdaA => P(4)(691),lamdaB => P(4)(755),s => s(4)(371),lamdaOut => P(3)(755));
U_G4756: entity G port map(lamdaA => P(4)(692),lamdaB => P(4)(756),s => s(4)(372),lamdaOut => P(3)(756));
U_G4757: entity G port map(lamdaA => P(4)(693),lamdaB => P(4)(757),s => s(4)(373),lamdaOut => P(3)(757));
U_G4758: entity G port map(lamdaA => P(4)(694),lamdaB => P(4)(758),s => s(4)(374),lamdaOut => P(3)(758));
U_G4759: entity G port map(lamdaA => P(4)(695),lamdaB => P(4)(759),s => s(4)(375),lamdaOut => P(3)(759));
U_G4760: entity G port map(lamdaA => P(4)(696),lamdaB => P(4)(760),s => s(4)(376),lamdaOut => P(3)(760));
U_G4761: entity G port map(lamdaA => P(4)(697),lamdaB => P(4)(761),s => s(4)(377),lamdaOut => P(3)(761));
U_G4762: entity G port map(lamdaA => P(4)(698),lamdaB => P(4)(762),s => s(4)(378),lamdaOut => P(3)(762));
U_G4763: entity G port map(lamdaA => P(4)(699),lamdaB => P(4)(763),s => s(4)(379),lamdaOut => P(3)(763));
U_G4764: entity G port map(lamdaA => P(4)(700),lamdaB => P(4)(764),s => s(4)(380),lamdaOut => P(3)(764));
U_G4765: entity G port map(lamdaA => P(4)(701),lamdaB => P(4)(765),s => s(4)(381),lamdaOut => P(3)(765));
U_G4766: entity G port map(lamdaA => P(4)(702),lamdaB => P(4)(766),s => s(4)(382),lamdaOut => P(3)(766));
U_G4767: entity G port map(lamdaA => P(4)(703),lamdaB => P(4)(767),s => s(4)(383),lamdaOut => P(3)(767));
U_F4768: entity F port map(lamdaA => P(4)(768),lamdaB => P(4)(832),lamdaOut => P(3)(768));
U_F4769: entity F port map(lamdaA => P(4)(769),lamdaB => P(4)(833),lamdaOut => P(3)(769));
U_F4770: entity F port map(lamdaA => P(4)(770),lamdaB => P(4)(834),lamdaOut => P(3)(770));
U_F4771: entity F port map(lamdaA => P(4)(771),lamdaB => P(4)(835),lamdaOut => P(3)(771));
U_F4772: entity F port map(lamdaA => P(4)(772),lamdaB => P(4)(836),lamdaOut => P(3)(772));
U_F4773: entity F port map(lamdaA => P(4)(773),lamdaB => P(4)(837),lamdaOut => P(3)(773));
U_F4774: entity F port map(lamdaA => P(4)(774),lamdaB => P(4)(838),lamdaOut => P(3)(774));
U_F4775: entity F port map(lamdaA => P(4)(775),lamdaB => P(4)(839),lamdaOut => P(3)(775));
U_F4776: entity F port map(lamdaA => P(4)(776),lamdaB => P(4)(840),lamdaOut => P(3)(776));
U_F4777: entity F port map(lamdaA => P(4)(777),lamdaB => P(4)(841),lamdaOut => P(3)(777));
U_F4778: entity F port map(lamdaA => P(4)(778),lamdaB => P(4)(842),lamdaOut => P(3)(778));
U_F4779: entity F port map(lamdaA => P(4)(779),lamdaB => P(4)(843),lamdaOut => P(3)(779));
U_F4780: entity F port map(lamdaA => P(4)(780),lamdaB => P(4)(844),lamdaOut => P(3)(780));
U_F4781: entity F port map(lamdaA => P(4)(781),lamdaB => P(4)(845),lamdaOut => P(3)(781));
U_F4782: entity F port map(lamdaA => P(4)(782),lamdaB => P(4)(846),lamdaOut => P(3)(782));
U_F4783: entity F port map(lamdaA => P(4)(783),lamdaB => P(4)(847),lamdaOut => P(3)(783));
U_F4784: entity F port map(lamdaA => P(4)(784),lamdaB => P(4)(848),lamdaOut => P(3)(784));
U_F4785: entity F port map(lamdaA => P(4)(785),lamdaB => P(4)(849),lamdaOut => P(3)(785));
U_F4786: entity F port map(lamdaA => P(4)(786),lamdaB => P(4)(850),lamdaOut => P(3)(786));
U_F4787: entity F port map(lamdaA => P(4)(787),lamdaB => P(4)(851),lamdaOut => P(3)(787));
U_F4788: entity F port map(lamdaA => P(4)(788),lamdaB => P(4)(852),lamdaOut => P(3)(788));
U_F4789: entity F port map(lamdaA => P(4)(789),lamdaB => P(4)(853),lamdaOut => P(3)(789));
U_F4790: entity F port map(lamdaA => P(4)(790),lamdaB => P(4)(854),lamdaOut => P(3)(790));
U_F4791: entity F port map(lamdaA => P(4)(791),lamdaB => P(4)(855),lamdaOut => P(3)(791));
U_F4792: entity F port map(lamdaA => P(4)(792),lamdaB => P(4)(856),lamdaOut => P(3)(792));
U_F4793: entity F port map(lamdaA => P(4)(793),lamdaB => P(4)(857),lamdaOut => P(3)(793));
U_F4794: entity F port map(lamdaA => P(4)(794),lamdaB => P(4)(858),lamdaOut => P(3)(794));
U_F4795: entity F port map(lamdaA => P(4)(795),lamdaB => P(4)(859),lamdaOut => P(3)(795));
U_F4796: entity F port map(lamdaA => P(4)(796),lamdaB => P(4)(860),lamdaOut => P(3)(796));
U_F4797: entity F port map(lamdaA => P(4)(797),lamdaB => P(4)(861),lamdaOut => P(3)(797));
U_F4798: entity F port map(lamdaA => P(4)(798),lamdaB => P(4)(862),lamdaOut => P(3)(798));
U_F4799: entity F port map(lamdaA => P(4)(799),lamdaB => P(4)(863),lamdaOut => P(3)(799));
U_F4800: entity F port map(lamdaA => P(4)(800),lamdaB => P(4)(864),lamdaOut => P(3)(800));
U_F4801: entity F port map(lamdaA => P(4)(801),lamdaB => P(4)(865),lamdaOut => P(3)(801));
U_F4802: entity F port map(lamdaA => P(4)(802),lamdaB => P(4)(866),lamdaOut => P(3)(802));
U_F4803: entity F port map(lamdaA => P(4)(803),lamdaB => P(4)(867),lamdaOut => P(3)(803));
U_F4804: entity F port map(lamdaA => P(4)(804),lamdaB => P(4)(868),lamdaOut => P(3)(804));
U_F4805: entity F port map(lamdaA => P(4)(805),lamdaB => P(4)(869),lamdaOut => P(3)(805));
U_F4806: entity F port map(lamdaA => P(4)(806),lamdaB => P(4)(870),lamdaOut => P(3)(806));
U_F4807: entity F port map(lamdaA => P(4)(807),lamdaB => P(4)(871),lamdaOut => P(3)(807));
U_F4808: entity F port map(lamdaA => P(4)(808),lamdaB => P(4)(872),lamdaOut => P(3)(808));
U_F4809: entity F port map(lamdaA => P(4)(809),lamdaB => P(4)(873),lamdaOut => P(3)(809));
U_F4810: entity F port map(lamdaA => P(4)(810),lamdaB => P(4)(874),lamdaOut => P(3)(810));
U_F4811: entity F port map(lamdaA => P(4)(811),lamdaB => P(4)(875),lamdaOut => P(3)(811));
U_F4812: entity F port map(lamdaA => P(4)(812),lamdaB => P(4)(876),lamdaOut => P(3)(812));
U_F4813: entity F port map(lamdaA => P(4)(813),lamdaB => P(4)(877),lamdaOut => P(3)(813));
U_F4814: entity F port map(lamdaA => P(4)(814),lamdaB => P(4)(878),lamdaOut => P(3)(814));
U_F4815: entity F port map(lamdaA => P(4)(815),lamdaB => P(4)(879),lamdaOut => P(3)(815));
U_F4816: entity F port map(lamdaA => P(4)(816),lamdaB => P(4)(880),lamdaOut => P(3)(816));
U_F4817: entity F port map(lamdaA => P(4)(817),lamdaB => P(4)(881),lamdaOut => P(3)(817));
U_F4818: entity F port map(lamdaA => P(4)(818),lamdaB => P(4)(882),lamdaOut => P(3)(818));
U_F4819: entity F port map(lamdaA => P(4)(819),lamdaB => P(4)(883),lamdaOut => P(3)(819));
U_F4820: entity F port map(lamdaA => P(4)(820),lamdaB => P(4)(884),lamdaOut => P(3)(820));
U_F4821: entity F port map(lamdaA => P(4)(821),lamdaB => P(4)(885),lamdaOut => P(3)(821));
U_F4822: entity F port map(lamdaA => P(4)(822),lamdaB => P(4)(886),lamdaOut => P(3)(822));
U_F4823: entity F port map(lamdaA => P(4)(823),lamdaB => P(4)(887),lamdaOut => P(3)(823));
U_F4824: entity F port map(lamdaA => P(4)(824),lamdaB => P(4)(888),lamdaOut => P(3)(824));
U_F4825: entity F port map(lamdaA => P(4)(825),lamdaB => P(4)(889),lamdaOut => P(3)(825));
U_F4826: entity F port map(lamdaA => P(4)(826),lamdaB => P(4)(890),lamdaOut => P(3)(826));
U_F4827: entity F port map(lamdaA => P(4)(827),lamdaB => P(4)(891),lamdaOut => P(3)(827));
U_F4828: entity F port map(lamdaA => P(4)(828),lamdaB => P(4)(892),lamdaOut => P(3)(828));
U_F4829: entity F port map(lamdaA => P(4)(829),lamdaB => P(4)(893),lamdaOut => P(3)(829));
U_F4830: entity F port map(lamdaA => P(4)(830),lamdaB => P(4)(894),lamdaOut => P(3)(830));
U_F4831: entity F port map(lamdaA => P(4)(831),lamdaB => P(4)(895),lamdaOut => P(3)(831));
U_G4832: entity G port map(lamdaA => P(4)(768),lamdaB => P(4)(832),s => s(4)(384),lamdaOut => P(3)(832));
U_G4833: entity G port map(lamdaA => P(4)(769),lamdaB => P(4)(833),s => s(4)(385),lamdaOut => P(3)(833));
U_G4834: entity G port map(lamdaA => P(4)(770),lamdaB => P(4)(834),s => s(4)(386),lamdaOut => P(3)(834));
U_G4835: entity G port map(lamdaA => P(4)(771),lamdaB => P(4)(835),s => s(4)(387),lamdaOut => P(3)(835));
U_G4836: entity G port map(lamdaA => P(4)(772),lamdaB => P(4)(836),s => s(4)(388),lamdaOut => P(3)(836));
U_G4837: entity G port map(lamdaA => P(4)(773),lamdaB => P(4)(837),s => s(4)(389),lamdaOut => P(3)(837));
U_G4838: entity G port map(lamdaA => P(4)(774),lamdaB => P(4)(838),s => s(4)(390),lamdaOut => P(3)(838));
U_G4839: entity G port map(lamdaA => P(4)(775),lamdaB => P(4)(839),s => s(4)(391),lamdaOut => P(3)(839));
U_G4840: entity G port map(lamdaA => P(4)(776),lamdaB => P(4)(840),s => s(4)(392),lamdaOut => P(3)(840));
U_G4841: entity G port map(lamdaA => P(4)(777),lamdaB => P(4)(841),s => s(4)(393),lamdaOut => P(3)(841));
U_G4842: entity G port map(lamdaA => P(4)(778),lamdaB => P(4)(842),s => s(4)(394),lamdaOut => P(3)(842));
U_G4843: entity G port map(lamdaA => P(4)(779),lamdaB => P(4)(843),s => s(4)(395),lamdaOut => P(3)(843));
U_G4844: entity G port map(lamdaA => P(4)(780),lamdaB => P(4)(844),s => s(4)(396),lamdaOut => P(3)(844));
U_G4845: entity G port map(lamdaA => P(4)(781),lamdaB => P(4)(845),s => s(4)(397),lamdaOut => P(3)(845));
U_G4846: entity G port map(lamdaA => P(4)(782),lamdaB => P(4)(846),s => s(4)(398),lamdaOut => P(3)(846));
U_G4847: entity G port map(lamdaA => P(4)(783),lamdaB => P(4)(847),s => s(4)(399),lamdaOut => P(3)(847));
U_G4848: entity G port map(lamdaA => P(4)(784),lamdaB => P(4)(848),s => s(4)(400),lamdaOut => P(3)(848));
U_G4849: entity G port map(lamdaA => P(4)(785),lamdaB => P(4)(849),s => s(4)(401),lamdaOut => P(3)(849));
U_G4850: entity G port map(lamdaA => P(4)(786),lamdaB => P(4)(850),s => s(4)(402),lamdaOut => P(3)(850));
U_G4851: entity G port map(lamdaA => P(4)(787),lamdaB => P(4)(851),s => s(4)(403),lamdaOut => P(3)(851));
U_G4852: entity G port map(lamdaA => P(4)(788),lamdaB => P(4)(852),s => s(4)(404),lamdaOut => P(3)(852));
U_G4853: entity G port map(lamdaA => P(4)(789),lamdaB => P(4)(853),s => s(4)(405),lamdaOut => P(3)(853));
U_G4854: entity G port map(lamdaA => P(4)(790),lamdaB => P(4)(854),s => s(4)(406),lamdaOut => P(3)(854));
U_G4855: entity G port map(lamdaA => P(4)(791),lamdaB => P(4)(855),s => s(4)(407),lamdaOut => P(3)(855));
U_G4856: entity G port map(lamdaA => P(4)(792),lamdaB => P(4)(856),s => s(4)(408),lamdaOut => P(3)(856));
U_G4857: entity G port map(lamdaA => P(4)(793),lamdaB => P(4)(857),s => s(4)(409),lamdaOut => P(3)(857));
U_G4858: entity G port map(lamdaA => P(4)(794),lamdaB => P(4)(858),s => s(4)(410),lamdaOut => P(3)(858));
U_G4859: entity G port map(lamdaA => P(4)(795),lamdaB => P(4)(859),s => s(4)(411),lamdaOut => P(3)(859));
U_G4860: entity G port map(lamdaA => P(4)(796),lamdaB => P(4)(860),s => s(4)(412),lamdaOut => P(3)(860));
U_G4861: entity G port map(lamdaA => P(4)(797),lamdaB => P(4)(861),s => s(4)(413),lamdaOut => P(3)(861));
U_G4862: entity G port map(lamdaA => P(4)(798),lamdaB => P(4)(862),s => s(4)(414),lamdaOut => P(3)(862));
U_G4863: entity G port map(lamdaA => P(4)(799),lamdaB => P(4)(863),s => s(4)(415),lamdaOut => P(3)(863));
U_G4864: entity G port map(lamdaA => P(4)(800),lamdaB => P(4)(864),s => s(4)(416),lamdaOut => P(3)(864));
U_G4865: entity G port map(lamdaA => P(4)(801),lamdaB => P(4)(865),s => s(4)(417),lamdaOut => P(3)(865));
U_G4866: entity G port map(lamdaA => P(4)(802),lamdaB => P(4)(866),s => s(4)(418),lamdaOut => P(3)(866));
U_G4867: entity G port map(lamdaA => P(4)(803),lamdaB => P(4)(867),s => s(4)(419),lamdaOut => P(3)(867));
U_G4868: entity G port map(lamdaA => P(4)(804),lamdaB => P(4)(868),s => s(4)(420),lamdaOut => P(3)(868));
U_G4869: entity G port map(lamdaA => P(4)(805),lamdaB => P(4)(869),s => s(4)(421),lamdaOut => P(3)(869));
U_G4870: entity G port map(lamdaA => P(4)(806),lamdaB => P(4)(870),s => s(4)(422),lamdaOut => P(3)(870));
U_G4871: entity G port map(lamdaA => P(4)(807),lamdaB => P(4)(871),s => s(4)(423),lamdaOut => P(3)(871));
U_G4872: entity G port map(lamdaA => P(4)(808),lamdaB => P(4)(872),s => s(4)(424),lamdaOut => P(3)(872));
U_G4873: entity G port map(lamdaA => P(4)(809),lamdaB => P(4)(873),s => s(4)(425),lamdaOut => P(3)(873));
U_G4874: entity G port map(lamdaA => P(4)(810),lamdaB => P(4)(874),s => s(4)(426),lamdaOut => P(3)(874));
U_G4875: entity G port map(lamdaA => P(4)(811),lamdaB => P(4)(875),s => s(4)(427),lamdaOut => P(3)(875));
U_G4876: entity G port map(lamdaA => P(4)(812),lamdaB => P(4)(876),s => s(4)(428),lamdaOut => P(3)(876));
U_G4877: entity G port map(lamdaA => P(4)(813),lamdaB => P(4)(877),s => s(4)(429),lamdaOut => P(3)(877));
U_G4878: entity G port map(lamdaA => P(4)(814),lamdaB => P(4)(878),s => s(4)(430),lamdaOut => P(3)(878));
U_G4879: entity G port map(lamdaA => P(4)(815),lamdaB => P(4)(879),s => s(4)(431),lamdaOut => P(3)(879));
U_G4880: entity G port map(lamdaA => P(4)(816),lamdaB => P(4)(880),s => s(4)(432),lamdaOut => P(3)(880));
U_G4881: entity G port map(lamdaA => P(4)(817),lamdaB => P(4)(881),s => s(4)(433),lamdaOut => P(3)(881));
U_G4882: entity G port map(lamdaA => P(4)(818),lamdaB => P(4)(882),s => s(4)(434),lamdaOut => P(3)(882));
U_G4883: entity G port map(lamdaA => P(4)(819),lamdaB => P(4)(883),s => s(4)(435),lamdaOut => P(3)(883));
U_G4884: entity G port map(lamdaA => P(4)(820),lamdaB => P(4)(884),s => s(4)(436),lamdaOut => P(3)(884));
U_G4885: entity G port map(lamdaA => P(4)(821),lamdaB => P(4)(885),s => s(4)(437),lamdaOut => P(3)(885));
U_G4886: entity G port map(lamdaA => P(4)(822),lamdaB => P(4)(886),s => s(4)(438),lamdaOut => P(3)(886));
U_G4887: entity G port map(lamdaA => P(4)(823),lamdaB => P(4)(887),s => s(4)(439),lamdaOut => P(3)(887));
U_G4888: entity G port map(lamdaA => P(4)(824),lamdaB => P(4)(888),s => s(4)(440),lamdaOut => P(3)(888));
U_G4889: entity G port map(lamdaA => P(4)(825),lamdaB => P(4)(889),s => s(4)(441),lamdaOut => P(3)(889));
U_G4890: entity G port map(lamdaA => P(4)(826),lamdaB => P(4)(890),s => s(4)(442),lamdaOut => P(3)(890));
U_G4891: entity G port map(lamdaA => P(4)(827),lamdaB => P(4)(891),s => s(4)(443),lamdaOut => P(3)(891));
U_G4892: entity G port map(lamdaA => P(4)(828),lamdaB => P(4)(892),s => s(4)(444),lamdaOut => P(3)(892));
U_G4893: entity G port map(lamdaA => P(4)(829),lamdaB => P(4)(893),s => s(4)(445),lamdaOut => P(3)(893));
U_G4894: entity G port map(lamdaA => P(4)(830),lamdaB => P(4)(894),s => s(4)(446),lamdaOut => P(3)(894));
U_G4895: entity G port map(lamdaA => P(4)(831),lamdaB => P(4)(895),s => s(4)(447),lamdaOut => P(3)(895));
U_F4896: entity F port map(lamdaA => P(4)(896),lamdaB => P(4)(960),lamdaOut => P(3)(896));
U_F4897: entity F port map(lamdaA => P(4)(897),lamdaB => P(4)(961),lamdaOut => P(3)(897));
U_F4898: entity F port map(lamdaA => P(4)(898),lamdaB => P(4)(962),lamdaOut => P(3)(898));
U_F4899: entity F port map(lamdaA => P(4)(899),lamdaB => P(4)(963),lamdaOut => P(3)(899));
U_F4900: entity F port map(lamdaA => P(4)(900),lamdaB => P(4)(964),lamdaOut => P(3)(900));
U_F4901: entity F port map(lamdaA => P(4)(901),lamdaB => P(4)(965),lamdaOut => P(3)(901));
U_F4902: entity F port map(lamdaA => P(4)(902),lamdaB => P(4)(966),lamdaOut => P(3)(902));
U_F4903: entity F port map(lamdaA => P(4)(903),lamdaB => P(4)(967),lamdaOut => P(3)(903));
U_F4904: entity F port map(lamdaA => P(4)(904),lamdaB => P(4)(968),lamdaOut => P(3)(904));
U_F4905: entity F port map(lamdaA => P(4)(905),lamdaB => P(4)(969),lamdaOut => P(3)(905));
U_F4906: entity F port map(lamdaA => P(4)(906),lamdaB => P(4)(970),lamdaOut => P(3)(906));
U_F4907: entity F port map(lamdaA => P(4)(907),lamdaB => P(4)(971),lamdaOut => P(3)(907));
U_F4908: entity F port map(lamdaA => P(4)(908),lamdaB => P(4)(972),lamdaOut => P(3)(908));
U_F4909: entity F port map(lamdaA => P(4)(909),lamdaB => P(4)(973),lamdaOut => P(3)(909));
U_F4910: entity F port map(lamdaA => P(4)(910),lamdaB => P(4)(974),lamdaOut => P(3)(910));
U_F4911: entity F port map(lamdaA => P(4)(911),lamdaB => P(4)(975),lamdaOut => P(3)(911));
U_F4912: entity F port map(lamdaA => P(4)(912),lamdaB => P(4)(976),lamdaOut => P(3)(912));
U_F4913: entity F port map(lamdaA => P(4)(913),lamdaB => P(4)(977),lamdaOut => P(3)(913));
U_F4914: entity F port map(lamdaA => P(4)(914),lamdaB => P(4)(978),lamdaOut => P(3)(914));
U_F4915: entity F port map(lamdaA => P(4)(915),lamdaB => P(4)(979),lamdaOut => P(3)(915));
U_F4916: entity F port map(lamdaA => P(4)(916),lamdaB => P(4)(980),lamdaOut => P(3)(916));
U_F4917: entity F port map(lamdaA => P(4)(917),lamdaB => P(4)(981),lamdaOut => P(3)(917));
U_F4918: entity F port map(lamdaA => P(4)(918),lamdaB => P(4)(982),lamdaOut => P(3)(918));
U_F4919: entity F port map(lamdaA => P(4)(919),lamdaB => P(4)(983),lamdaOut => P(3)(919));
U_F4920: entity F port map(lamdaA => P(4)(920),lamdaB => P(4)(984),lamdaOut => P(3)(920));
U_F4921: entity F port map(lamdaA => P(4)(921),lamdaB => P(4)(985),lamdaOut => P(3)(921));
U_F4922: entity F port map(lamdaA => P(4)(922),lamdaB => P(4)(986),lamdaOut => P(3)(922));
U_F4923: entity F port map(lamdaA => P(4)(923),lamdaB => P(4)(987),lamdaOut => P(3)(923));
U_F4924: entity F port map(lamdaA => P(4)(924),lamdaB => P(4)(988),lamdaOut => P(3)(924));
U_F4925: entity F port map(lamdaA => P(4)(925),lamdaB => P(4)(989),lamdaOut => P(3)(925));
U_F4926: entity F port map(lamdaA => P(4)(926),lamdaB => P(4)(990),lamdaOut => P(3)(926));
U_F4927: entity F port map(lamdaA => P(4)(927),lamdaB => P(4)(991),lamdaOut => P(3)(927));
U_F4928: entity F port map(lamdaA => P(4)(928),lamdaB => P(4)(992),lamdaOut => P(3)(928));
U_F4929: entity F port map(lamdaA => P(4)(929),lamdaB => P(4)(993),lamdaOut => P(3)(929));
U_F4930: entity F port map(lamdaA => P(4)(930),lamdaB => P(4)(994),lamdaOut => P(3)(930));
U_F4931: entity F port map(lamdaA => P(4)(931),lamdaB => P(4)(995),lamdaOut => P(3)(931));
U_F4932: entity F port map(lamdaA => P(4)(932),lamdaB => P(4)(996),lamdaOut => P(3)(932));
U_F4933: entity F port map(lamdaA => P(4)(933),lamdaB => P(4)(997),lamdaOut => P(3)(933));
U_F4934: entity F port map(lamdaA => P(4)(934),lamdaB => P(4)(998),lamdaOut => P(3)(934));
U_F4935: entity F port map(lamdaA => P(4)(935),lamdaB => P(4)(999),lamdaOut => P(3)(935));
U_F4936: entity F port map(lamdaA => P(4)(936),lamdaB => P(4)(1000),lamdaOut => P(3)(936));
U_F4937: entity F port map(lamdaA => P(4)(937),lamdaB => P(4)(1001),lamdaOut => P(3)(937));
U_F4938: entity F port map(lamdaA => P(4)(938),lamdaB => P(4)(1002),lamdaOut => P(3)(938));
U_F4939: entity F port map(lamdaA => P(4)(939),lamdaB => P(4)(1003),lamdaOut => P(3)(939));
U_F4940: entity F port map(lamdaA => P(4)(940),lamdaB => P(4)(1004),lamdaOut => P(3)(940));
U_F4941: entity F port map(lamdaA => P(4)(941),lamdaB => P(4)(1005),lamdaOut => P(3)(941));
U_F4942: entity F port map(lamdaA => P(4)(942),lamdaB => P(4)(1006),lamdaOut => P(3)(942));
U_F4943: entity F port map(lamdaA => P(4)(943),lamdaB => P(4)(1007),lamdaOut => P(3)(943));
U_F4944: entity F port map(lamdaA => P(4)(944),lamdaB => P(4)(1008),lamdaOut => P(3)(944));
U_F4945: entity F port map(lamdaA => P(4)(945),lamdaB => P(4)(1009),lamdaOut => P(3)(945));
U_F4946: entity F port map(lamdaA => P(4)(946),lamdaB => P(4)(1010),lamdaOut => P(3)(946));
U_F4947: entity F port map(lamdaA => P(4)(947),lamdaB => P(4)(1011),lamdaOut => P(3)(947));
U_F4948: entity F port map(lamdaA => P(4)(948),lamdaB => P(4)(1012),lamdaOut => P(3)(948));
U_F4949: entity F port map(lamdaA => P(4)(949),lamdaB => P(4)(1013),lamdaOut => P(3)(949));
U_F4950: entity F port map(lamdaA => P(4)(950),lamdaB => P(4)(1014),lamdaOut => P(3)(950));
U_F4951: entity F port map(lamdaA => P(4)(951),lamdaB => P(4)(1015),lamdaOut => P(3)(951));
U_F4952: entity F port map(lamdaA => P(4)(952),lamdaB => P(4)(1016),lamdaOut => P(3)(952));
U_F4953: entity F port map(lamdaA => P(4)(953),lamdaB => P(4)(1017),lamdaOut => P(3)(953));
U_F4954: entity F port map(lamdaA => P(4)(954),lamdaB => P(4)(1018),lamdaOut => P(3)(954));
U_F4955: entity F port map(lamdaA => P(4)(955),lamdaB => P(4)(1019),lamdaOut => P(3)(955));
U_F4956: entity F port map(lamdaA => P(4)(956),lamdaB => P(4)(1020),lamdaOut => P(3)(956));
U_F4957: entity F port map(lamdaA => P(4)(957),lamdaB => P(4)(1021),lamdaOut => P(3)(957));
U_F4958: entity F port map(lamdaA => P(4)(958),lamdaB => P(4)(1022),lamdaOut => P(3)(958));
U_F4959: entity F port map(lamdaA => P(4)(959),lamdaB => P(4)(1023),lamdaOut => P(3)(959));
U_G4960: entity G port map(lamdaA => P(4)(896),lamdaB => P(4)(960),s => s(4)(448),lamdaOut => P(3)(960));
U_G4961: entity G port map(lamdaA => P(4)(897),lamdaB => P(4)(961),s => s(4)(449),lamdaOut => P(3)(961));
U_G4962: entity G port map(lamdaA => P(4)(898),lamdaB => P(4)(962),s => s(4)(450),lamdaOut => P(3)(962));
U_G4963: entity G port map(lamdaA => P(4)(899),lamdaB => P(4)(963),s => s(4)(451),lamdaOut => P(3)(963));
U_G4964: entity G port map(lamdaA => P(4)(900),lamdaB => P(4)(964),s => s(4)(452),lamdaOut => P(3)(964));
U_G4965: entity G port map(lamdaA => P(4)(901),lamdaB => P(4)(965),s => s(4)(453),lamdaOut => P(3)(965));
U_G4966: entity G port map(lamdaA => P(4)(902),lamdaB => P(4)(966),s => s(4)(454),lamdaOut => P(3)(966));
U_G4967: entity G port map(lamdaA => P(4)(903),lamdaB => P(4)(967),s => s(4)(455),lamdaOut => P(3)(967));
U_G4968: entity G port map(lamdaA => P(4)(904),lamdaB => P(4)(968),s => s(4)(456),lamdaOut => P(3)(968));
U_G4969: entity G port map(lamdaA => P(4)(905),lamdaB => P(4)(969),s => s(4)(457),lamdaOut => P(3)(969));
U_G4970: entity G port map(lamdaA => P(4)(906),lamdaB => P(4)(970),s => s(4)(458),lamdaOut => P(3)(970));
U_G4971: entity G port map(lamdaA => P(4)(907),lamdaB => P(4)(971),s => s(4)(459),lamdaOut => P(3)(971));
U_G4972: entity G port map(lamdaA => P(4)(908),lamdaB => P(4)(972),s => s(4)(460),lamdaOut => P(3)(972));
U_G4973: entity G port map(lamdaA => P(4)(909),lamdaB => P(4)(973),s => s(4)(461),lamdaOut => P(3)(973));
U_G4974: entity G port map(lamdaA => P(4)(910),lamdaB => P(4)(974),s => s(4)(462),lamdaOut => P(3)(974));
U_G4975: entity G port map(lamdaA => P(4)(911),lamdaB => P(4)(975),s => s(4)(463),lamdaOut => P(3)(975));
U_G4976: entity G port map(lamdaA => P(4)(912),lamdaB => P(4)(976),s => s(4)(464),lamdaOut => P(3)(976));
U_G4977: entity G port map(lamdaA => P(4)(913),lamdaB => P(4)(977),s => s(4)(465),lamdaOut => P(3)(977));
U_G4978: entity G port map(lamdaA => P(4)(914),lamdaB => P(4)(978),s => s(4)(466),lamdaOut => P(3)(978));
U_G4979: entity G port map(lamdaA => P(4)(915),lamdaB => P(4)(979),s => s(4)(467),lamdaOut => P(3)(979));
U_G4980: entity G port map(lamdaA => P(4)(916),lamdaB => P(4)(980),s => s(4)(468),lamdaOut => P(3)(980));
U_G4981: entity G port map(lamdaA => P(4)(917),lamdaB => P(4)(981),s => s(4)(469),lamdaOut => P(3)(981));
U_G4982: entity G port map(lamdaA => P(4)(918),lamdaB => P(4)(982),s => s(4)(470),lamdaOut => P(3)(982));
U_G4983: entity G port map(lamdaA => P(4)(919),lamdaB => P(4)(983),s => s(4)(471),lamdaOut => P(3)(983));
U_G4984: entity G port map(lamdaA => P(4)(920),lamdaB => P(4)(984),s => s(4)(472),lamdaOut => P(3)(984));
U_G4985: entity G port map(lamdaA => P(4)(921),lamdaB => P(4)(985),s => s(4)(473),lamdaOut => P(3)(985));
U_G4986: entity G port map(lamdaA => P(4)(922),lamdaB => P(4)(986),s => s(4)(474),lamdaOut => P(3)(986));
U_G4987: entity G port map(lamdaA => P(4)(923),lamdaB => P(4)(987),s => s(4)(475),lamdaOut => P(3)(987));
U_G4988: entity G port map(lamdaA => P(4)(924),lamdaB => P(4)(988),s => s(4)(476),lamdaOut => P(3)(988));
U_G4989: entity G port map(lamdaA => P(4)(925),lamdaB => P(4)(989),s => s(4)(477),lamdaOut => P(3)(989));
U_G4990: entity G port map(lamdaA => P(4)(926),lamdaB => P(4)(990),s => s(4)(478),lamdaOut => P(3)(990));
U_G4991: entity G port map(lamdaA => P(4)(927),lamdaB => P(4)(991),s => s(4)(479),lamdaOut => P(3)(991));
U_G4992: entity G port map(lamdaA => P(4)(928),lamdaB => P(4)(992),s => s(4)(480),lamdaOut => P(3)(992));
U_G4993: entity G port map(lamdaA => P(4)(929),lamdaB => P(4)(993),s => s(4)(481),lamdaOut => P(3)(993));
U_G4994: entity G port map(lamdaA => P(4)(930),lamdaB => P(4)(994),s => s(4)(482),lamdaOut => P(3)(994));
U_G4995: entity G port map(lamdaA => P(4)(931),lamdaB => P(4)(995),s => s(4)(483),lamdaOut => P(3)(995));
U_G4996: entity G port map(lamdaA => P(4)(932),lamdaB => P(4)(996),s => s(4)(484),lamdaOut => P(3)(996));
U_G4997: entity G port map(lamdaA => P(4)(933),lamdaB => P(4)(997),s => s(4)(485),lamdaOut => P(3)(997));
U_G4998: entity G port map(lamdaA => P(4)(934),lamdaB => P(4)(998),s => s(4)(486),lamdaOut => P(3)(998));
U_G4999: entity G port map(lamdaA => P(4)(935),lamdaB => P(4)(999),s => s(4)(487),lamdaOut => P(3)(999));
U_G41000: entity G port map(lamdaA => P(4)(936),lamdaB => P(4)(1000),s => s(4)(488),lamdaOut => P(3)(1000));
U_G41001: entity G port map(lamdaA => P(4)(937),lamdaB => P(4)(1001),s => s(4)(489),lamdaOut => P(3)(1001));
U_G41002: entity G port map(lamdaA => P(4)(938),lamdaB => P(4)(1002),s => s(4)(490),lamdaOut => P(3)(1002));
U_G41003: entity G port map(lamdaA => P(4)(939),lamdaB => P(4)(1003),s => s(4)(491),lamdaOut => P(3)(1003));
U_G41004: entity G port map(lamdaA => P(4)(940),lamdaB => P(4)(1004),s => s(4)(492),lamdaOut => P(3)(1004));
U_G41005: entity G port map(lamdaA => P(4)(941),lamdaB => P(4)(1005),s => s(4)(493),lamdaOut => P(3)(1005));
U_G41006: entity G port map(lamdaA => P(4)(942),lamdaB => P(4)(1006),s => s(4)(494),lamdaOut => P(3)(1006));
U_G41007: entity G port map(lamdaA => P(4)(943),lamdaB => P(4)(1007),s => s(4)(495),lamdaOut => P(3)(1007));
U_G41008: entity G port map(lamdaA => P(4)(944),lamdaB => P(4)(1008),s => s(4)(496),lamdaOut => P(3)(1008));
U_G41009: entity G port map(lamdaA => P(4)(945),lamdaB => P(4)(1009),s => s(4)(497),lamdaOut => P(3)(1009));
U_G41010: entity G port map(lamdaA => P(4)(946),lamdaB => P(4)(1010),s => s(4)(498),lamdaOut => P(3)(1010));
U_G41011: entity G port map(lamdaA => P(4)(947),lamdaB => P(4)(1011),s => s(4)(499),lamdaOut => P(3)(1011));
U_G41012: entity G port map(lamdaA => P(4)(948),lamdaB => P(4)(1012),s => s(4)(500),lamdaOut => P(3)(1012));
U_G41013: entity G port map(lamdaA => P(4)(949),lamdaB => P(4)(1013),s => s(4)(501),lamdaOut => P(3)(1013));
U_G41014: entity G port map(lamdaA => P(4)(950),lamdaB => P(4)(1014),s => s(4)(502),lamdaOut => P(3)(1014));
U_G41015: entity G port map(lamdaA => P(4)(951),lamdaB => P(4)(1015),s => s(4)(503),lamdaOut => P(3)(1015));
U_G41016: entity G port map(lamdaA => P(4)(952),lamdaB => P(4)(1016),s => s(4)(504),lamdaOut => P(3)(1016));
U_G41017: entity G port map(lamdaA => P(4)(953),lamdaB => P(4)(1017),s => s(4)(505),lamdaOut => P(3)(1017));
U_G41018: entity G port map(lamdaA => P(4)(954),lamdaB => P(4)(1018),s => s(4)(506),lamdaOut => P(3)(1018));
U_G41019: entity G port map(lamdaA => P(4)(955),lamdaB => P(4)(1019),s => s(4)(507),lamdaOut => P(3)(1019));
U_G41020: entity G port map(lamdaA => P(4)(956),lamdaB => P(4)(1020),s => s(4)(508),lamdaOut => P(3)(1020));
U_G41021: entity G port map(lamdaA => P(4)(957),lamdaB => P(4)(1021),s => s(4)(509),lamdaOut => P(3)(1021));
U_G41022: entity G port map(lamdaA => P(4)(958),lamdaB => P(4)(1022),s => s(4)(510),lamdaOut => P(3)(1022));
U_G41023: entity G port map(lamdaA => P(4)(959),lamdaB => P(4)(1023),s => s(4)(511),lamdaOut => P(3)(1023));
-- STAGE 2
U_F30: entity F port map(lamdaA => P(3)(0),lamdaB => P(3)(128),lamdaOut => P(2)(0));
U_F31: entity F port map(lamdaA => P(3)(1),lamdaB => P(3)(129),lamdaOut => P(2)(1));
U_F32: entity F port map(lamdaA => P(3)(2),lamdaB => P(3)(130),lamdaOut => P(2)(2));
U_F33: entity F port map(lamdaA => P(3)(3),lamdaB => P(3)(131),lamdaOut => P(2)(3));
U_F34: entity F port map(lamdaA => P(3)(4),lamdaB => P(3)(132),lamdaOut => P(2)(4));
U_F35: entity F port map(lamdaA => P(3)(5),lamdaB => P(3)(133),lamdaOut => P(2)(5));
U_F36: entity F port map(lamdaA => P(3)(6),lamdaB => P(3)(134),lamdaOut => P(2)(6));
U_F37: entity F port map(lamdaA => P(3)(7),lamdaB => P(3)(135),lamdaOut => P(2)(7));
U_F38: entity F port map(lamdaA => P(3)(8),lamdaB => P(3)(136),lamdaOut => P(2)(8));
U_F39: entity F port map(lamdaA => P(3)(9),lamdaB => P(3)(137),lamdaOut => P(2)(9));
U_F310: entity F port map(lamdaA => P(3)(10),lamdaB => P(3)(138),lamdaOut => P(2)(10));
U_F311: entity F port map(lamdaA => P(3)(11),lamdaB => P(3)(139),lamdaOut => P(2)(11));
U_F312: entity F port map(lamdaA => P(3)(12),lamdaB => P(3)(140),lamdaOut => P(2)(12));
U_F313: entity F port map(lamdaA => P(3)(13),lamdaB => P(3)(141),lamdaOut => P(2)(13));
U_F314: entity F port map(lamdaA => P(3)(14),lamdaB => P(3)(142),lamdaOut => P(2)(14));
U_F315: entity F port map(lamdaA => P(3)(15),lamdaB => P(3)(143),lamdaOut => P(2)(15));
U_F316: entity F port map(lamdaA => P(3)(16),lamdaB => P(3)(144),lamdaOut => P(2)(16));
U_F317: entity F port map(lamdaA => P(3)(17),lamdaB => P(3)(145),lamdaOut => P(2)(17));
U_F318: entity F port map(lamdaA => P(3)(18),lamdaB => P(3)(146),lamdaOut => P(2)(18));
U_F319: entity F port map(lamdaA => P(3)(19),lamdaB => P(3)(147),lamdaOut => P(2)(19));
U_F320: entity F port map(lamdaA => P(3)(20),lamdaB => P(3)(148),lamdaOut => P(2)(20));
U_F321: entity F port map(lamdaA => P(3)(21),lamdaB => P(3)(149),lamdaOut => P(2)(21));
U_F322: entity F port map(lamdaA => P(3)(22),lamdaB => P(3)(150),lamdaOut => P(2)(22));
U_F323: entity F port map(lamdaA => P(3)(23),lamdaB => P(3)(151),lamdaOut => P(2)(23));
U_F324: entity F port map(lamdaA => P(3)(24),lamdaB => P(3)(152),lamdaOut => P(2)(24));
U_F325: entity F port map(lamdaA => P(3)(25),lamdaB => P(3)(153),lamdaOut => P(2)(25));
U_F326: entity F port map(lamdaA => P(3)(26),lamdaB => P(3)(154),lamdaOut => P(2)(26));
U_F327: entity F port map(lamdaA => P(3)(27),lamdaB => P(3)(155),lamdaOut => P(2)(27));
U_F328: entity F port map(lamdaA => P(3)(28),lamdaB => P(3)(156),lamdaOut => P(2)(28));
U_F329: entity F port map(lamdaA => P(3)(29),lamdaB => P(3)(157),lamdaOut => P(2)(29));
U_F330: entity F port map(lamdaA => P(3)(30),lamdaB => P(3)(158),lamdaOut => P(2)(30));
U_F331: entity F port map(lamdaA => P(3)(31),lamdaB => P(3)(159),lamdaOut => P(2)(31));
U_F332: entity F port map(lamdaA => P(3)(32),lamdaB => P(3)(160),lamdaOut => P(2)(32));
U_F333: entity F port map(lamdaA => P(3)(33),lamdaB => P(3)(161),lamdaOut => P(2)(33));
U_F334: entity F port map(lamdaA => P(3)(34),lamdaB => P(3)(162),lamdaOut => P(2)(34));
U_F335: entity F port map(lamdaA => P(3)(35),lamdaB => P(3)(163),lamdaOut => P(2)(35));
U_F336: entity F port map(lamdaA => P(3)(36),lamdaB => P(3)(164),lamdaOut => P(2)(36));
U_F337: entity F port map(lamdaA => P(3)(37),lamdaB => P(3)(165),lamdaOut => P(2)(37));
U_F338: entity F port map(lamdaA => P(3)(38),lamdaB => P(3)(166),lamdaOut => P(2)(38));
U_F339: entity F port map(lamdaA => P(3)(39),lamdaB => P(3)(167),lamdaOut => P(2)(39));
U_F340: entity F port map(lamdaA => P(3)(40),lamdaB => P(3)(168),lamdaOut => P(2)(40));
U_F341: entity F port map(lamdaA => P(3)(41),lamdaB => P(3)(169),lamdaOut => P(2)(41));
U_F342: entity F port map(lamdaA => P(3)(42),lamdaB => P(3)(170),lamdaOut => P(2)(42));
U_F343: entity F port map(lamdaA => P(3)(43),lamdaB => P(3)(171),lamdaOut => P(2)(43));
U_F344: entity F port map(lamdaA => P(3)(44),lamdaB => P(3)(172),lamdaOut => P(2)(44));
U_F345: entity F port map(lamdaA => P(3)(45),lamdaB => P(3)(173),lamdaOut => P(2)(45));
U_F346: entity F port map(lamdaA => P(3)(46),lamdaB => P(3)(174),lamdaOut => P(2)(46));
U_F347: entity F port map(lamdaA => P(3)(47),lamdaB => P(3)(175),lamdaOut => P(2)(47));
U_F348: entity F port map(lamdaA => P(3)(48),lamdaB => P(3)(176),lamdaOut => P(2)(48));
U_F349: entity F port map(lamdaA => P(3)(49),lamdaB => P(3)(177),lamdaOut => P(2)(49));
U_F350: entity F port map(lamdaA => P(3)(50),lamdaB => P(3)(178),lamdaOut => P(2)(50));
U_F351: entity F port map(lamdaA => P(3)(51),lamdaB => P(3)(179),lamdaOut => P(2)(51));
U_F352: entity F port map(lamdaA => P(3)(52),lamdaB => P(3)(180),lamdaOut => P(2)(52));
U_F353: entity F port map(lamdaA => P(3)(53),lamdaB => P(3)(181),lamdaOut => P(2)(53));
U_F354: entity F port map(lamdaA => P(3)(54),lamdaB => P(3)(182),lamdaOut => P(2)(54));
U_F355: entity F port map(lamdaA => P(3)(55),lamdaB => P(3)(183),lamdaOut => P(2)(55));
U_F356: entity F port map(lamdaA => P(3)(56),lamdaB => P(3)(184),lamdaOut => P(2)(56));
U_F357: entity F port map(lamdaA => P(3)(57),lamdaB => P(3)(185),lamdaOut => P(2)(57));
U_F358: entity F port map(lamdaA => P(3)(58),lamdaB => P(3)(186),lamdaOut => P(2)(58));
U_F359: entity F port map(lamdaA => P(3)(59),lamdaB => P(3)(187),lamdaOut => P(2)(59));
U_F360: entity F port map(lamdaA => P(3)(60),lamdaB => P(3)(188),lamdaOut => P(2)(60));
U_F361: entity F port map(lamdaA => P(3)(61),lamdaB => P(3)(189),lamdaOut => P(2)(61));
U_F362: entity F port map(lamdaA => P(3)(62),lamdaB => P(3)(190),lamdaOut => P(2)(62));
U_F363: entity F port map(lamdaA => P(3)(63),lamdaB => P(3)(191),lamdaOut => P(2)(63));
U_F364: entity F port map(lamdaA => P(3)(64),lamdaB => P(3)(192),lamdaOut => P(2)(64));
U_F365: entity F port map(lamdaA => P(3)(65),lamdaB => P(3)(193),lamdaOut => P(2)(65));
U_F366: entity F port map(lamdaA => P(3)(66),lamdaB => P(3)(194),lamdaOut => P(2)(66));
U_F367: entity F port map(lamdaA => P(3)(67),lamdaB => P(3)(195),lamdaOut => P(2)(67));
U_F368: entity F port map(lamdaA => P(3)(68),lamdaB => P(3)(196),lamdaOut => P(2)(68));
U_F369: entity F port map(lamdaA => P(3)(69),lamdaB => P(3)(197),lamdaOut => P(2)(69));
U_F370: entity F port map(lamdaA => P(3)(70),lamdaB => P(3)(198),lamdaOut => P(2)(70));
U_F371: entity F port map(lamdaA => P(3)(71),lamdaB => P(3)(199),lamdaOut => P(2)(71));
U_F372: entity F port map(lamdaA => P(3)(72),lamdaB => P(3)(200),lamdaOut => P(2)(72));
U_F373: entity F port map(lamdaA => P(3)(73),lamdaB => P(3)(201),lamdaOut => P(2)(73));
U_F374: entity F port map(lamdaA => P(3)(74),lamdaB => P(3)(202),lamdaOut => P(2)(74));
U_F375: entity F port map(lamdaA => P(3)(75),lamdaB => P(3)(203),lamdaOut => P(2)(75));
U_F376: entity F port map(lamdaA => P(3)(76),lamdaB => P(3)(204),lamdaOut => P(2)(76));
U_F377: entity F port map(lamdaA => P(3)(77),lamdaB => P(3)(205),lamdaOut => P(2)(77));
U_F378: entity F port map(lamdaA => P(3)(78),lamdaB => P(3)(206),lamdaOut => P(2)(78));
U_F379: entity F port map(lamdaA => P(3)(79),lamdaB => P(3)(207),lamdaOut => P(2)(79));
U_F380: entity F port map(lamdaA => P(3)(80),lamdaB => P(3)(208),lamdaOut => P(2)(80));
U_F381: entity F port map(lamdaA => P(3)(81),lamdaB => P(3)(209),lamdaOut => P(2)(81));
U_F382: entity F port map(lamdaA => P(3)(82),lamdaB => P(3)(210),lamdaOut => P(2)(82));
U_F383: entity F port map(lamdaA => P(3)(83),lamdaB => P(3)(211),lamdaOut => P(2)(83));
U_F384: entity F port map(lamdaA => P(3)(84),lamdaB => P(3)(212),lamdaOut => P(2)(84));
U_F385: entity F port map(lamdaA => P(3)(85),lamdaB => P(3)(213),lamdaOut => P(2)(85));
U_F386: entity F port map(lamdaA => P(3)(86),lamdaB => P(3)(214),lamdaOut => P(2)(86));
U_F387: entity F port map(lamdaA => P(3)(87),lamdaB => P(3)(215),lamdaOut => P(2)(87));
U_F388: entity F port map(lamdaA => P(3)(88),lamdaB => P(3)(216),lamdaOut => P(2)(88));
U_F389: entity F port map(lamdaA => P(3)(89),lamdaB => P(3)(217),lamdaOut => P(2)(89));
U_F390: entity F port map(lamdaA => P(3)(90),lamdaB => P(3)(218),lamdaOut => P(2)(90));
U_F391: entity F port map(lamdaA => P(3)(91),lamdaB => P(3)(219),lamdaOut => P(2)(91));
U_F392: entity F port map(lamdaA => P(3)(92),lamdaB => P(3)(220),lamdaOut => P(2)(92));
U_F393: entity F port map(lamdaA => P(3)(93),lamdaB => P(3)(221),lamdaOut => P(2)(93));
U_F394: entity F port map(lamdaA => P(3)(94),lamdaB => P(3)(222),lamdaOut => P(2)(94));
U_F395: entity F port map(lamdaA => P(3)(95),lamdaB => P(3)(223),lamdaOut => P(2)(95));
U_F396: entity F port map(lamdaA => P(3)(96),lamdaB => P(3)(224),lamdaOut => P(2)(96));
U_F397: entity F port map(lamdaA => P(3)(97),lamdaB => P(3)(225),lamdaOut => P(2)(97));
U_F398: entity F port map(lamdaA => P(3)(98),lamdaB => P(3)(226),lamdaOut => P(2)(98));
U_F399: entity F port map(lamdaA => P(3)(99),lamdaB => P(3)(227),lamdaOut => P(2)(99));
U_F3100: entity F port map(lamdaA => P(3)(100),lamdaB => P(3)(228),lamdaOut => P(2)(100));
U_F3101: entity F port map(lamdaA => P(3)(101),lamdaB => P(3)(229),lamdaOut => P(2)(101));
U_F3102: entity F port map(lamdaA => P(3)(102),lamdaB => P(3)(230),lamdaOut => P(2)(102));
U_F3103: entity F port map(lamdaA => P(3)(103),lamdaB => P(3)(231),lamdaOut => P(2)(103));
U_F3104: entity F port map(lamdaA => P(3)(104),lamdaB => P(3)(232),lamdaOut => P(2)(104));
U_F3105: entity F port map(lamdaA => P(3)(105),lamdaB => P(3)(233),lamdaOut => P(2)(105));
U_F3106: entity F port map(lamdaA => P(3)(106),lamdaB => P(3)(234),lamdaOut => P(2)(106));
U_F3107: entity F port map(lamdaA => P(3)(107),lamdaB => P(3)(235),lamdaOut => P(2)(107));
U_F3108: entity F port map(lamdaA => P(3)(108),lamdaB => P(3)(236),lamdaOut => P(2)(108));
U_F3109: entity F port map(lamdaA => P(3)(109),lamdaB => P(3)(237),lamdaOut => P(2)(109));
U_F3110: entity F port map(lamdaA => P(3)(110),lamdaB => P(3)(238),lamdaOut => P(2)(110));
U_F3111: entity F port map(lamdaA => P(3)(111),lamdaB => P(3)(239),lamdaOut => P(2)(111));
U_F3112: entity F port map(lamdaA => P(3)(112),lamdaB => P(3)(240),lamdaOut => P(2)(112));
U_F3113: entity F port map(lamdaA => P(3)(113),lamdaB => P(3)(241),lamdaOut => P(2)(113));
U_F3114: entity F port map(lamdaA => P(3)(114),lamdaB => P(3)(242),lamdaOut => P(2)(114));
U_F3115: entity F port map(lamdaA => P(3)(115),lamdaB => P(3)(243),lamdaOut => P(2)(115));
U_F3116: entity F port map(lamdaA => P(3)(116),lamdaB => P(3)(244),lamdaOut => P(2)(116));
U_F3117: entity F port map(lamdaA => P(3)(117),lamdaB => P(3)(245),lamdaOut => P(2)(117));
U_F3118: entity F port map(lamdaA => P(3)(118),lamdaB => P(3)(246),lamdaOut => P(2)(118));
U_F3119: entity F port map(lamdaA => P(3)(119),lamdaB => P(3)(247),lamdaOut => P(2)(119));
U_F3120: entity F port map(lamdaA => P(3)(120),lamdaB => P(3)(248),lamdaOut => P(2)(120));
U_F3121: entity F port map(lamdaA => P(3)(121),lamdaB => P(3)(249),lamdaOut => P(2)(121));
U_F3122: entity F port map(lamdaA => P(3)(122),lamdaB => P(3)(250),lamdaOut => P(2)(122));
U_F3123: entity F port map(lamdaA => P(3)(123),lamdaB => P(3)(251),lamdaOut => P(2)(123));
U_F3124: entity F port map(lamdaA => P(3)(124),lamdaB => P(3)(252),lamdaOut => P(2)(124));
U_F3125: entity F port map(lamdaA => P(3)(125),lamdaB => P(3)(253),lamdaOut => P(2)(125));
U_F3126: entity F port map(lamdaA => P(3)(126),lamdaB => P(3)(254),lamdaOut => P(2)(126));
U_F3127: entity F port map(lamdaA => P(3)(127),lamdaB => P(3)(255),lamdaOut => P(2)(127));
U_G3128: entity G port map(lamdaA => P(3)(0),lamdaB => P(3)(128),s => s(3)(0),lamdaOut => P(2)(128));
U_G3129: entity G port map(lamdaA => P(3)(1),lamdaB => P(3)(129),s => s(3)(1),lamdaOut => P(2)(129));
U_G3130: entity G port map(lamdaA => P(3)(2),lamdaB => P(3)(130),s => s(3)(2),lamdaOut => P(2)(130));
U_G3131: entity G port map(lamdaA => P(3)(3),lamdaB => P(3)(131),s => s(3)(3),lamdaOut => P(2)(131));
U_G3132: entity G port map(lamdaA => P(3)(4),lamdaB => P(3)(132),s => s(3)(4),lamdaOut => P(2)(132));
U_G3133: entity G port map(lamdaA => P(3)(5),lamdaB => P(3)(133),s => s(3)(5),lamdaOut => P(2)(133));
U_G3134: entity G port map(lamdaA => P(3)(6),lamdaB => P(3)(134),s => s(3)(6),lamdaOut => P(2)(134));
U_G3135: entity G port map(lamdaA => P(3)(7),lamdaB => P(3)(135),s => s(3)(7),lamdaOut => P(2)(135));
U_G3136: entity G port map(lamdaA => P(3)(8),lamdaB => P(3)(136),s => s(3)(8),lamdaOut => P(2)(136));
U_G3137: entity G port map(lamdaA => P(3)(9),lamdaB => P(3)(137),s => s(3)(9),lamdaOut => P(2)(137));
U_G3138: entity G port map(lamdaA => P(3)(10),lamdaB => P(3)(138),s => s(3)(10),lamdaOut => P(2)(138));
U_G3139: entity G port map(lamdaA => P(3)(11),lamdaB => P(3)(139),s => s(3)(11),lamdaOut => P(2)(139));
U_G3140: entity G port map(lamdaA => P(3)(12),lamdaB => P(3)(140),s => s(3)(12),lamdaOut => P(2)(140));
U_G3141: entity G port map(lamdaA => P(3)(13),lamdaB => P(3)(141),s => s(3)(13),lamdaOut => P(2)(141));
U_G3142: entity G port map(lamdaA => P(3)(14),lamdaB => P(3)(142),s => s(3)(14),lamdaOut => P(2)(142));
U_G3143: entity G port map(lamdaA => P(3)(15),lamdaB => P(3)(143),s => s(3)(15),lamdaOut => P(2)(143));
U_G3144: entity G port map(lamdaA => P(3)(16),lamdaB => P(3)(144),s => s(3)(16),lamdaOut => P(2)(144));
U_G3145: entity G port map(lamdaA => P(3)(17),lamdaB => P(3)(145),s => s(3)(17),lamdaOut => P(2)(145));
U_G3146: entity G port map(lamdaA => P(3)(18),lamdaB => P(3)(146),s => s(3)(18),lamdaOut => P(2)(146));
U_G3147: entity G port map(lamdaA => P(3)(19),lamdaB => P(3)(147),s => s(3)(19),lamdaOut => P(2)(147));
U_G3148: entity G port map(lamdaA => P(3)(20),lamdaB => P(3)(148),s => s(3)(20),lamdaOut => P(2)(148));
U_G3149: entity G port map(lamdaA => P(3)(21),lamdaB => P(3)(149),s => s(3)(21),lamdaOut => P(2)(149));
U_G3150: entity G port map(lamdaA => P(3)(22),lamdaB => P(3)(150),s => s(3)(22),lamdaOut => P(2)(150));
U_G3151: entity G port map(lamdaA => P(3)(23),lamdaB => P(3)(151),s => s(3)(23),lamdaOut => P(2)(151));
U_G3152: entity G port map(lamdaA => P(3)(24),lamdaB => P(3)(152),s => s(3)(24),lamdaOut => P(2)(152));
U_G3153: entity G port map(lamdaA => P(3)(25),lamdaB => P(3)(153),s => s(3)(25),lamdaOut => P(2)(153));
U_G3154: entity G port map(lamdaA => P(3)(26),lamdaB => P(3)(154),s => s(3)(26),lamdaOut => P(2)(154));
U_G3155: entity G port map(lamdaA => P(3)(27),lamdaB => P(3)(155),s => s(3)(27),lamdaOut => P(2)(155));
U_G3156: entity G port map(lamdaA => P(3)(28),lamdaB => P(3)(156),s => s(3)(28),lamdaOut => P(2)(156));
U_G3157: entity G port map(lamdaA => P(3)(29),lamdaB => P(3)(157),s => s(3)(29),lamdaOut => P(2)(157));
U_G3158: entity G port map(lamdaA => P(3)(30),lamdaB => P(3)(158),s => s(3)(30),lamdaOut => P(2)(158));
U_G3159: entity G port map(lamdaA => P(3)(31),lamdaB => P(3)(159),s => s(3)(31),lamdaOut => P(2)(159));
U_G3160: entity G port map(lamdaA => P(3)(32),lamdaB => P(3)(160),s => s(3)(32),lamdaOut => P(2)(160));
U_G3161: entity G port map(lamdaA => P(3)(33),lamdaB => P(3)(161),s => s(3)(33),lamdaOut => P(2)(161));
U_G3162: entity G port map(lamdaA => P(3)(34),lamdaB => P(3)(162),s => s(3)(34),lamdaOut => P(2)(162));
U_G3163: entity G port map(lamdaA => P(3)(35),lamdaB => P(3)(163),s => s(3)(35),lamdaOut => P(2)(163));
U_G3164: entity G port map(lamdaA => P(3)(36),lamdaB => P(3)(164),s => s(3)(36),lamdaOut => P(2)(164));
U_G3165: entity G port map(lamdaA => P(3)(37),lamdaB => P(3)(165),s => s(3)(37),lamdaOut => P(2)(165));
U_G3166: entity G port map(lamdaA => P(3)(38),lamdaB => P(3)(166),s => s(3)(38),lamdaOut => P(2)(166));
U_G3167: entity G port map(lamdaA => P(3)(39),lamdaB => P(3)(167),s => s(3)(39),lamdaOut => P(2)(167));
U_G3168: entity G port map(lamdaA => P(3)(40),lamdaB => P(3)(168),s => s(3)(40),lamdaOut => P(2)(168));
U_G3169: entity G port map(lamdaA => P(3)(41),lamdaB => P(3)(169),s => s(3)(41),lamdaOut => P(2)(169));
U_G3170: entity G port map(lamdaA => P(3)(42),lamdaB => P(3)(170),s => s(3)(42),lamdaOut => P(2)(170));
U_G3171: entity G port map(lamdaA => P(3)(43),lamdaB => P(3)(171),s => s(3)(43),lamdaOut => P(2)(171));
U_G3172: entity G port map(lamdaA => P(3)(44),lamdaB => P(3)(172),s => s(3)(44),lamdaOut => P(2)(172));
U_G3173: entity G port map(lamdaA => P(3)(45),lamdaB => P(3)(173),s => s(3)(45),lamdaOut => P(2)(173));
U_G3174: entity G port map(lamdaA => P(3)(46),lamdaB => P(3)(174),s => s(3)(46),lamdaOut => P(2)(174));
U_G3175: entity G port map(lamdaA => P(3)(47),lamdaB => P(3)(175),s => s(3)(47),lamdaOut => P(2)(175));
U_G3176: entity G port map(lamdaA => P(3)(48),lamdaB => P(3)(176),s => s(3)(48),lamdaOut => P(2)(176));
U_G3177: entity G port map(lamdaA => P(3)(49),lamdaB => P(3)(177),s => s(3)(49),lamdaOut => P(2)(177));
U_G3178: entity G port map(lamdaA => P(3)(50),lamdaB => P(3)(178),s => s(3)(50),lamdaOut => P(2)(178));
U_G3179: entity G port map(lamdaA => P(3)(51),lamdaB => P(3)(179),s => s(3)(51),lamdaOut => P(2)(179));
U_G3180: entity G port map(lamdaA => P(3)(52),lamdaB => P(3)(180),s => s(3)(52),lamdaOut => P(2)(180));
U_G3181: entity G port map(lamdaA => P(3)(53),lamdaB => P(3)(181),s => s(3)(53),lamdaOut => P(2)(181));
U_G3182: entity G port map(lamdaA => P(3)(54),lamdaB => P(3)(182),s => s(3)(54),lamdaOut => P(2)(182));
U_G3183: entity G port map(lamdaA => P(3)(55),lamdaB => P(3)(183),s => s(3)(55),lamdaOut => P(2)(183));
U_G3184: entity G port map(lamdaA => P(3)(56),lamdaB => P(3)(184),s => s(3)(56),lamdaOut => P(2)(184));
U_G3185: entity G port map(lamdaA => P(3)(57),lamdaB => P(3)(185),s => s(3)(57),lamdaOut => P(2)(185));
U_G3186: entity G port map(lamdaA => P(3)(58),lamdaB => P(3)(186),s => s(3)(58),lamdaOut => P(2)(186));
U_G3187: entity G port map(lamdaA => P(3)(59),lamdaB => P(3)(187),s => s(3)(59),lamdaOut => P(2)(187));
U_G3188: entity G port map(lamdaA => P(3)(60),lamdaB => P(3)(188),s => s(3)(60),lamdaOut => P(2)(188));
U_G3189: entity G port map(lamdaA => P(3)(61),lamdaB => P(3)(189),s => s(3)(61),lamdaOut => P(2)(189));
U_G3190: entity G port map(lamdaA => P(3)(62),lamdaB => P(3)(190),s => s(3)(62),lamdaOut => P(2)(190));
U_G3191: entity G port map(lamdaA => P(3)(63),lamdaB => P(3)(191),s => s(3)(63),lamdaOut => P(2)(191));
U_G3192: entity G port map(lamdaA => P(3)(64),lamdaB => P(3)(192),s => s(3)(64),lamdaOut => P(2)(192));
U_G3193: entity G port map(lamdaA => P(3)(65),lamdaB => P(3)(193),s => s(3)(65),lamdaOut => P(2)(193));
U_G3194: entity G port map(lamdaA => P(3)(66),lamdaB => P(3)(194),s => s(3)(66),lamdaOut => P(2)(194));
U_G3195: entity G port map(lamdaA => P(3)(67),lamdaB => P(3)(195),s => s(3)(67),lamdaOut => P(2)(195));
U_G3196: entity G port map(lamdaA => P(3)(68),lamdaB => P(3)(196),s => s(3)(68),lamdaOut => P(2)(196));
U_G3197: entity G port map(lamdaA => P(3)(69),lamdaB => P(3)(197),s => s(3)(69),lamdaOut => P(2)(197));
U_G3198: entity G port map(lamdaA => P(3)(70),lamdaB => P(3)(198),s => s(3)(70),lamdaOut => P(2)(198));
U_G3199: entity G port map(lamdaA => P(3)(71),lamdaB => P(3)(199),s => s(3)(71),lamdaOut => P(2)(199));
U_G3200: entity G port map(lamdaA => P(3)(72),lamdaB => P(3)(200),s => s(3)(72),lamdaOut => P(2)(200));
U_G3201: entity G port map(lamdaA => P(3)(73),lamdaB => P(3)(201),s => s(3)(73),lamdaOut => P(2)(201));
U_G3202: entity G port map(lamdaA => P(3)(74),lamdaB => P(3)(202),s => s(3)(74),lamdaOut => P(2)(202));
U_G3203: entity G port map(lamdaA => P(3)(75),lamdaB => P(3)(203),s => s(3)(75),lamdaOut => P(2)(203));
U_G3204: entity G port map(lamdaA => P(3)(76),lamdaB => P(3)(204),s => s(3)(76),lamdaOut => P(2)(204));
U_G3205: entity G port map(lamdaA => P(3)(77),lamdaB => P(3)(205),s => s(3)(77),lamdaOut => P(2)(205));
U_G3206: entity G port map(lamdaA => P(3)(78),lamdaB => P(3)(206),s => s(3)(78),lamdaOut => P(2)(206));
U_G3207: entity G port map(lamdaA => P(3)(79),lamdaB => P(3)(207),s => s(3)(79),lamdaOut => P(2)(207));
U_G3208: entity G port map(lamdaA => P(3)(80),lamdaB => P(3)(208),s => s(3)(80),lamdaOut => P(2)(208));
U_G3209: entity G port map(lamdaA => P(3)(81),lamdaB => P(3)(209),s => s(3)(81),lamdaOut => P(2)(209));
U_G3210: entity G port map(lamdaA => P(3)(82),lamdaB => P(3)(210),s => s(3)(82),lamdaOut => P(2)(210));
U_G3211: entity G port map(lamdaA => P(3)(83),lamdaB => P(3)(211),s => s(3)(83),lamdaOut => P(2)(211));
U_G3212: entity G port map(lamdaA => P(3)(84),lamdaB => P(3)(212),s => s(3)(84),lamdaOut => P(2)(212));
U_G3213: entity G port map(lamdaA => P(3)(85),lamdaB => P(3)(213),s => s(3)(85),lamdaOut => P(2)(213));
U_G3214: entity G port map(lamdaA => P(3)(86),lamdaB => P(3)(214),s => s(3)(86),lamdaOut => P(2)(214));
U_G3215: entity G port map(lamdaA => P(3)(87),lamdaB => P(3)(215),s => s(3)(87),lamdaOut => P(2)(215));
U_G3216: entity G port map(lamdaA => P(3)(88),lamdaB => P(3)(216),s => s(3)(88),lamdaOut => P(2)(216));
U_G3217: entity G port map(lamdaA => P(3)(89),lamdaB => P(3)(217),s => s(3)(89),lamdaOut => P(2)(217));
U_G3218: entity G port map(lamdaA => P(3)(90),lamdaB => P(3)(218),s => s(3)(90),lamdaOut => P(2)(218));
U_G3219: entity G port map(lamdaA => P(3)(91),lamdaB => P(3)(219),s => s(3)(91),lamdaOut => P(2)(219));
U_G3220: entity G port map(lamdaA => P(3)(92),lamdaB => P(3)(220),s => s(3)(92),lamdaOut => P(2)(220));
U_G3221: entity G port map(lamdaA => P(3)(93),lamdaB => P(3)(221),s => s(3)(93),lamdaOut => P(2)(221));
U_G3222: entity G port map(lamdaA => P(3)(94),lamdaB => P(3)(222),s => s(3)(94),lamdaOut => P(2)(222));
U_G3223: entity G port map(lamdaA => P(3)(95),lamdaB => P(3)(223),s => s(3)(95),lamdaOut => P(2)(223));
U_G3224: entity G port map(lamdaA => P(3)(96),lamdaB => P(3)(224),s => s(3)(96),lamdaOut => P(2)(224));
U_G3225: entity G port map(lamdaA => P(3)(97),lamdaB => P(3)(225),s => s(3)(97),lamdaOut => P(2)(225));
U_G3226: entity G port map(lamdaA => P(3)(98),lamdaB => P(3)(226),s => s(3)(98),lamdaOut => P(2)(226));
U_G3227: entity G port map(lamdaA => P(3)(99),lamdaB => P(3)(227),s => s(3)(99),lamdaOut => P(2)(227));
U_G3228: entity G port map(lamdaA => P(3)(100),lamdaB => P(3)(228),s => s(3)(100),lamdaOut => P(2)(228));
U_G3229: entity G port map(lamdaA => P(3)(101),lamdaB => P(3)(229),s => s(3)(101),lamdaOut => P(2)(229));
U_G3230: entity G port map(lamdaA => P(3)(102),lamdaB => P(3)(230),s => s(3)(102),lamdaOut => P(2)(230));
U_G3231: entity G port map(lamdaA => P(3)(103),lamdaB => P(3)(231),s => s(3)(103),lamdaOut => P(2)(231));
U_G3232: entity G port map(lamdaA => P(3)(104),lamdaB => P(3)(232),s => s(3)(104),lamdaOut => P(2)(232));
U_G3233: entity G port map(lamdaA => P(3)(105),lamdaB => P(3)(233),s => s(3)(105),lamdaOut => P(2)(233));
U_G3234: entity G port map(lamdaA => P(3)(106),lamdaB => P(3)(234),s => s(3)(106),lamdaOut => P(2)(234));
U_G3235: entity G port map(lamdaA => P(3)(107),lamdaB => P(3)(235),s => s(3)(107),lamdaOut => P(2)(235));
U_G3236: entity G port map(lamdaA => P(3)(108),lamdaB => P(3)(236),s => s(3)(108),lamdaOut => P(2)(236));
U_G3237: entity G port map(lamdaA => P(3)(109),lamdaB => P(3)(237),s => s(3)(109),lamdaOut => P(2)(237));
U_G3238: entity G port map(lamdaA => P(3)(110),lamdaB => P(3)(238),s => s(3)(110),lamdaOut => P(2)(238));
U_G3239: entity G port map(lamdaA => P(3)(111),lamdaB => P(3)(239),s => s(3)(111),lamdaOut => P(2)(239));
U_G3240: entity G port map(lamdaA => P(3)(112),lamdaB => P(3)(240),s => s(3)(112),lamdaOut => P(2)(240));
U_G3241: entity G port map(lamdaA => P(3)(113),lamdaB => P(3)(241),s => s(3)(113),lamdaOut => P(2)(241));
U_G3242: entity G port map(lamdaA => P(3)(114),lamdaB => P(3)(242),s => s(3)(114),lamdaOut => P(2)(242));
U_G3243: entity G port map(lamdaA => P(3)(115),lamdaB => P(3)(243),s => s(3)(115),lamdaOut => P(2)(243));
U_G3244: entity G port map(lamdaA => P(3)(116),lamdaB => P(3)(244),s => s(3)(116),lamdaOut => P(2)(244));
U_G3245: entity G port map(lamdaA => P(3)(117),lamdaB => P(3)(245),s => s(3)(117),lamdaOut => P(2)(245));
U_G3246: entity G port map(lamdaA => P(3)(118),lamdaB => P(3)(246),s => s(3)(118),lamdaOut => P(2)(246));
U_G3247: entity G port map(lamdaA => P(3)(119),lamdaB => P(3)(247),s => s(3)(119),lamdaOut => P(2)(247));
U_G3248: entity G port map(lamdaA => P(3)(120),lamdaB => P(3)(248),s => s(3)(120),lamdaOut => P(2)(248));
U_G3249: entity G port map(lamdaA => P(3)(121),lamdaB => P(3)(249),s => s(3)(121),lamdaOut => P(2)(249));
U_G3250: entity G port map(lamdaA => P(3)(122),lamdaB => P(3)(250),s => s(3)(122),lamdaOut => P(2)(250));
U_G3251: entity G port map(lamdaA => P(3)(123),lamdaB => P(3)(251),s => s(3)(123),lamdaOut => P(2)(251));
U_G3252: entity G port map(lamdaA => P(3)(124),lamdaB => P(3)(252),s => s(3)(124),lamdaOut => P(2)(252));
U_G3253: entity G port map(lamdaA => P(3)(125),lamdaB => P(3)(253),s => s(3)(125),lamdaOut => P(2)(253));
U_G3254: entity G port map(lamdaA => P(3)(126),lamdaB => P(3)(254),s => s(3)(126),lamdaOut => P(2)(254));
U_G3255: entity G port map(lamdaA => P(3)(127),lamdaB => P(3)(255),s => s(3)(127),lamdaOut => P(2)(255));
U_F3256: entity F port map(lamdaA => P(3)(256),lamdaB => P(3)(384),lamdaOut => P(2)(256));
U_F3257: entity F port map(lamdaA => P(3)(257),lamdaB => P(3)(385),lamdaOut => P(2)(257));
U_F3258: entity F port map(lamdaA => P(3)(258),lamdaB => P(3)(386),lamdaOut => P(2)(258));
U_F3259: entity F port map(lamdaA => P(3)(259),lamdaB => P(3)(387),lamdaOut => P(2)(259));
U_F3260: entity F port map(lamdaA => P(3)(260),lamdaB => P(3)(388),lamdaOut => P(2)(260));
U_F3261: entity F port map(lamdaA => P(3)(261),lamdaB => P(3)(389),lamdaOut => P(2)(261));
U_F3262: entity F port map(lamdaA => P(3)(262),lamdaB => P(3)(390),lamdaOut => P(2)(262));
U_F3263: entity F port map(lamdaA => P(3)(263),lamdaB => P(3)(391),lamdaOut => P(2)(263));
U_F3264: entity F port map(lamdaA => P(3)(264),lamdaB => P(3)(392),lamdaOut => P(2)(264));
U_F3265: entity F port map(lamdaA => P(3)(265),lamdaB => P(3)(393),lamdaOut => P(2)(265));
U_F3266: entity F port map(lamdaA => P(3)(266),lamdaB => P(3)(394),lamdaOut => P(2)(266));
U_F3267: entity F port map(lamdaA => P(3)(267),lamdaB => P(3)(395),lamdaOut => P(2)(267));
U_F3268: entity F port map(lamdaA => P(3)(268),lamdaB => P(3)(396),lamdaOut => P(2)(268));
U_F3269: entity F port map(lamdaA => P(3)(269),lamdaB => P(3)(397),lamdaOut => P(2)(269));
U_F3270: entity F port map(lamdaA => P(3)(270),lamdaB => P(3)(398),lamdaOut => P(2)(270));
U_F3271: entity F port map(lamdaA => P(3)(271),lamdaB => P(3)(399),lamdaOut => P(2)(271));
U_F3272: entity F port map(lamdaA => P(3)(272),lamdaB => P(3)(400),lamdaOut => P(2)(272));
U_F3273: entity F port map(lamdaA => P(3)(273),lamdaB => P(3)(401),lamdaOut => P(2)(273));
U_F3274: entity F port map(lamdaA => P(3)(274),lamdaB => P(3)(402),lamdaOut => P(2)(274));
U_F3275: entity F port map(lamdaA => P(3)(275),lamdaB => P(3)(403),lamdaOut => P(2)(275));
U_F3276: entity F port map(lamdaA => P(3)(276),lamdaB => P(3)(404),lamdaOut => P(2)(276));
U_F3277: entity F port map(lamdaA => P(3)(277),lamdaB => P(3)(405),lamdaOut => P(2)(277));
U_F3278: entity F port map(lamdaA => P(3)(278),lamdaB => P(3)(406),lamdaOut => P(2)(278));
U_F3279: entity F port map(lamdaA => P(3)(279),lamdaB => P(3)(407),lamdaOut => P(2)(279));
U_F3280: entity F port map(lamdaA => P(3)(280),lamdaB => P(3)(408),lamdaOut => P(2)(280));
U_F3281: entity F port map(lamdaA => P(3)(281),lamdaB => P(3)(409),lamdaOut => P(2)(281));
U_F3282: entity F port map(lamdaA => P(3)(282),lamdaB => P(3)(410),lamdaOut => P(2)(282));
U_F3283: entity F port map(lamdaA => P(3)(283),lamdaB => P(3)(411),lamdaOut => P(2)(283));
U_F3284: entity F port map(lamdaA => P(3)(284),lamdaB => P(3)(412),lamdaOut => P(2)(284));
U_F3285: entity F port map(lamdaA => P(3)(285),lamdaB => P(3)(413),lamdaOut => P(2)(285));
U_F3286: entity F port map(lamdaA => P(3)(286),lamdaB => P(3)(414),lamdaOut => P(2)(286));
U_F3287: entity F port map(lamdaA => P(3)(287),lamdaB => P(3)(415),lamdaOut => P(2)(287));
U_F3288: entity F port map(lamdaA => P(3)(288),lamdaB => P(3)(416),lamdaOut => P(2)(288));
U_F3289: entity F port map(lamdaA => P(3)(289),lamdaB => P(3)(417),lamdaOut => P(2)(289));
U_F3290: entity F port map(lamdaA => P(3)(290),lamdaB => P(3)(418),lamdaOut => P(2)(290));
U_F3291: entity F port map(lamdaA => P(3)(291),lamdaB => P(3)(419),lamdaOut => P(2)(291));
U_F3292: entity F port map(lamdaA => P(3)(292),lamdaB => P(3)(420),lamdaOut => P(2)(292));
U_F3293: entity F port map(lamdaA => P(3)(293),lamdaB => P(3)(421),lamdaOut => P(2)(293));
U_F3294: entity F port map(lamdaA => P(3)(294),lamdaB => P(3)(422),lamdaOut => P(2)(294));
U_F3295: entity F port map(lamdaA => P(3)(295),lamdaB => P(3)(423),lamdaOut => P(2)(295));
U_F3296: entity F port map(lamdaA => P(3)(296),lamdaB => P(3)(424),lamdaOut => P(2)(296));
U_F3297: entity F port map(lamdaA => P(3)(297),lamdaB => P(3)(425),lamdaOut => P(2)(297));
U_F3298: entity F port map(lamdaA => P(3)(298),lamdaB => P(3)(426),lamdaOut => P(2)(298));
U_F3299: entity F port map(lamdaA => P(3)(299),lamdaB => P(3)(427),lamdaOut => P(2)(299));
U_F3300: entity F port map(lamdaA => P(3)(300),lamdaB => P(3)(428),lamdaOut => P(2)(300));
U_F3301: entity F port map(lamdaA => P(3)(301),lamdaB => P(3)(429),lamdaOut => P(2)(301));
U_F3302: entity F port map(lamdaA => P(3)(302),lamdaB => P(3)(430),lamdaOut => P(2)(302));
U_F3303: entity F port map(lamdaA => P(3)(303),lamdaB => P(3)(431),lamdaOut => P(2)(303));
U_F3304: entity F port map(lamdaA => P(3)(304),lamdaB => P(3)(432),lamdaOut => P(2)(304));
U_F3305: entity F port map(lamdaA => P(3)(305),lamdaB => P(3)(433),lamdaOut => P(2)(305));
U_F3306: entity F port map(lamdaA => P(3)(306),lamdaB => P(3)(434),lamdaOut => P(2)(306));
U_F3307: entity F port map(lamdaA => P(3)(307),lamdaB => P(3)(435),lamdaOut => P(2)(307));
U_F3308: entity F port map(lamdaA => P(3)(308),lamdaB => P(3)(436),lamdaOut => P(2)(308));
U_F3309: entity F port map(lamdaA => P(3)(309),lamdaB => P(3)(437),lamdaOut => P(2)(309));
U_F3310: entity F port map(lamdaA => P(3)(310),lamdaB => P(3)(438),lamdaOut => P(2)(310));
U_F3311: entity F port map(lamdaA => P(3)(311),lamdaB => P(3)(439),lamdaOut => P(2)(311));
U_F3312: entity F port map(lamdaA => P(3)(312),lamdaB => P(3)(440),lamdaOut => P(2)(312));
U_F3313: entity F port map(lamdaA => P(3)(313),lamdaB => P(3)(441),lamdaOut => P(2)(313));
U_F3314: entity F port map(lamdaA => P(3)(314),lamdaB => P(3)(442),lamdaOut => P(2)(314));
U_F3315: entity F port map(lamdaA => P(3)(315),lamdaB => P(3)(443),lamdaOut => P(2)(315));
U_F3316: entity F port map(lamdaA => P(3)(316),lamdaB => P(3)(444),lamdaOut => P(2)(316));
U_F3317: entity F port map(lamdaA => P(3)(317),lamdaB => P(3)(445),lamdaOut => P(2)(317));
U_F3318: entity F port map(lamdaA => P(3)(318),lamdaB => P(3)(446),lamdaOut => P(2)(318));
U_F3319: entity F port map(lamdaA => P(3)(319),lamdaB => P(3)(447),lamdaOut => P(2)(319));
U_F3320: entity F port map(lamdaA => P(3)(320),lamdaB => P(3)(448),lamdaOut => P(2)(320));
U_F3321: entity F port map(lamdaA => P(3)(321),lamdaB => P(3)(449),lamdaOut => P(2)(321));
U_F3322: entity F port map(lamdaA => P(3)(322),lamdaB => P(3)(450),lamdaOut => P(2)(322));
U_F3323: entity F port map(lamdaA => P(3)(323),lamdaB => P(3)(451),lamdaOut => P(2)(323));
U_F3324: entity F port map(lamdaA => P(3)(324),lamdaB => P(3)(452),lamdaOut => P(2)(324));
U_F3325: entity F port map(lamdaA => P(3)(325),lamdaB => P(3)(453),lamdaOut => P(2)(325));
U_F3326: entity F port map(lamdaA => P(3)(326),lamdaB => P(3)(454),lamdaOut => P(2)(326));
U_F3327: entity F port map(lamdaA => P(3)(327),lamdaB => P(3)(455),lamdaOut => P(2)(327));
U_F3328: entity F port map(lamdaA => P(3)(328),lamdaB => P(3)(456),lamdaOut => P(2)(328));
U_F3329: entity F port map(lamdaA => P(3)(329),lamdaB => P(3)(457),lamdaOut => P(2)(329));
U_F3330: entity F port map(lamdaA => P(3)(330),lamdaB => P(3)(458),lamdaOut => P(2)(330));
U_F3331: entity F port map(lamdaA => P(3)(331),lamdaB => P(3)(459),lamdaOut => P(2)(331));
U_F3332: entity F port map(lamdaA => P(3)(332),lamdaB => P(3)(460),lamdaOut => P(2)(332));
U_F3333: entity F port map(lamdaA => P(3)(333),lamdaB => P(3)(461),lamdaOut => P(2)(333));
U_F3334: entity F port map(lamdaA => P(3)(334),lamdaB => P(3)(462),lamdaOut => P(2)(334));
U_F3335: entity F port map(lamdaA => P(3)(335),lamdaB => P(3)(463),lamdaOut => P(2)(335));
U_F3336: entity F port map(lamdaA => P(3)(336),lamdaB => P(3)(464),lamdaOut => P(2)(336));
U_F3337: entity F port map(lamdaA => P(3)(337),lamdaB => P(3)(465),lamdaOut => P(2)(337));
U_F3338: entity F port map(lamdaA => P(3)(338),lamdaB => P(3)(466),lamdaOut => P(2)(338));
U_F3339: entity F port map(lamdaA => P(3)(339),lamdaB => P(3)(467),lamdaOut => P(2)(339));
U_F3340: entity F port map(lamdaA => P(3)(340),lamdaB => P(3)(468),lamdaOut => P(2)(340));
U_F3341: entity F port map(lamdaA => P(3)(341),lamdaB => P(3)(469),lamdaOut => P(2)(341));
U_F3342: entity F port map(lamdaA => P(3)(342),lamdaB => P(3)(470),lamdaOut => P(2)(342));
U_F3343: entity F port map(lamdaA => P(3)(343),lamdaB => P(3)(471),lamdaOut => P(2)(343));
U_F3344: entity F port map(lamdaA => P(3)(344),lamdaB => P(3)(472),lamdaOut => P(2)(344));
U_F3345: entity F port map(lamdaA => P(3)(345),lamdaB => P(3)(473),lamdaOut => P(2)(345));
U_F3346: entity F port map(lamdaA => P(3)(346),lamdaB => P(3)(474),lamdaOut => P(2)(346));
U_F3347: entity F port map(lamdaA => P(3)(347),lamdaB => P(3)(475),lamdaOut => P(2)(347));
U_F3348: entity F port map(lamdaA => P(3)(348),lamdaB => P(3)(476),lamdaOut => P(2)(348));
U_F3349: entity F port map(lamdaA => P(3)(349),lamdaB => P(3)(477),lamdaOut => P(2)(349));
U_F3350: entity F port map(lamdaA => P(3)(350),lamdaB => P(3)(478),lamdaOut => P(2)(350));
U_F3351: entity F port map(lamdaA => P(3)(351),lamdaB => P(3)(479),lamdaOut => P(2)(351));
U_F3352: entity F port map(lamdaA => P(3)(352),lamdaB => P(3)(480),lamdaOut => P(2)(352));
U_F3353: entity F port map(lamdaA => P(3)(353),lamdaB => P(3)(481),lamdaOut => P(2)(353));
U_F3354: entity F port map(lamdaA => P(3)(354),lamdaB => P(3)(482),lamdaOut => P(2)(354));
U_F3355: entity F port map(lamdaA => P(3)(355),lamdaB => P(3)(483),lamdaOut => P(2)(355));
U_F3356: entity F port map(lamdaA => P(3)(356),lamdaB => P(3)(484),lamdaOut => P(2)(356));
U_F3357: entity F port map(lamdaA => P(3)(357),lamdaB => P(3)(485),lamdaOut => P(2)(357));
U_F3358: entity F port map(lamdaA => P(3)(358),lamdaB => P(3)(486),lamdaOut => P(2)(358));
U_F3359: entity F port map(lamdaA => P(3)(359),lamdaB => P(3)(487),lamdaOut => P(2)(359));
U_F3360: entity F port map(lamdaA => P(3)(360),lamdaB => P(3)(488),lamdaOut => P(2)(360));
U_F3361: entity F port map(lamdaA => P(3)(361),lamdaB => P(3)(489),lamdaOut => P(2)(361));
U_F3362: entity F port map(lamdaA => P(3)(362),lamdaB => P(3)(490),lamdaOut => P(2)(362));
U_F3363: entity F port map(lamdaA => P(3)(363),lamdaB => P(3)(491),lamdaOut => P(2)(363));
U_F3364: entity F port map(lamdaA => P(3)(364),lamdaB => P(3)(492),lamdaOut => P(2)(364));
U_F3365: entity F port map(lamdaA => P(3)(365),lamdaB => P(3)(493),lamdaOut => P(2)(365));
U_F3366: entity F port map(lamdaA => P(3)(366),lamdaB => P(3)(494),lamdaOut => P(2)(366));
U_F3367: entity F port map(lamdaA => P(3)(367),lamdaB => P(3)(495),lamdaOut => P(2)(367));
U_F3368: entity F port map(lamdaA => P(3)(368),lamdaB => P(3)(496),lamdaOut => P(2)(368));
U_F3369: entity F port map(lamdaA => P(3)(369),lamdaB => P(3)(497),lamdaOut => P(2)(369));
U_F3370: entity F port map(lamdaA => P(3)(370),lamdaB => P(3)(498),lamdaOut => P(2)(370));
U_F3371: entity F port map(lamdaA => P(3)(371),lamdaB => P(3)(499),lamdaOut => P(2)(371));
U_F3372: entity F port map(lamdaA => P(3)(372),lamdaB => P(3)(500),lamdaOut => P(2)(372));
U_F3373: entity F port map(lamdaA => P(3)(373),lamdaB => P(3)(501),lamdaOut => P(2)(373));
U_F3374: entity F port map(lamdaA => P(3)(374),lamdaB => P(3)(502),lamdaOut => P(2)(374));
U_F3375: entity F port map(lamdaA => P(3)(375),lamdaB => P(3)(503),lamdaOut => P(2)(375));
U_F3376: entity F port map(lamdaA => P(3)(376),lamdaB => P(3)(504),lamdaOut => P(2)(376));
U_F3377: entity F port map(lamdaA => P(3)(377),lamdaB => P(3)(505),lamdaOut => P(2)(377));
U_F3378: entity F port map(lamdaA => P(3)(378),lamdaB => P(3)(506),lamdaOut => P(2)(378));
U_F3379: entity F port map(lamdaA => P(3)(379),lamdaB => P(3)(507),lamdaOut => P(2)(379));
U_F3380: entity F port map(lamdaA => P(3)(380),lamdaB => P(3)(508),lamdaOut => P(2)(380));
U_F3381: entity F port map(lamdaA => P(3)(381),lamdaB => P(3)(509),lamdaOut => P(2)(381));
U_F3382: entity F port map(lamdaA => P(3)(382),lamdaB => P(3)(510),lamdaOut => P(2)(382));
U_F3383: entity F port map(lamdaA => P(3)(383),lamdaB => P(3)(511),lamdaOut => P(2)(383));
U_G3384: entity G port map(lamdaA => P(3)(256),lamdaB => P(3)(384),s => s(3)(128),lamdaOut => P(2)(384));
U_G3385: entity G port map(lamdaA => P(3)(257),lamdaB => P(3)(385),s => s(3)(129),lamdaOut => P(2)(385));
U_G3386: entity G port map(lamdaA => P(3)(258),lamdaB => P(3)(386),s => s(3)(130),lamdaOut => P(2)(386));
U_G3387: entity G port map(lamdaA => P(3)(259),lamdaB => P(3)(387),s => s(3)(131),lamdaOut => P(2)(387));
U_G3388: entity G port map(lamdaA => P(3)(260),lamdaB => P(3)(388),s => s(3)(132),lamdaOut => P(2)(388));
U_G3389: entity G port map(lamdaA => P(3)(261),lamdaB => P(3)(389),s => s(3)(133),lamdaOut => P(2)(389));
U_G3390: entity G port map(lamdaA => P(3)(262),lamdaB => P(3)(390),s => s(3)(134),lamdaOut => P(2)(390));
U_G3391: entity G port map(lamdaA => P(3)(263),lamdaB => P(3)(391),s => s(3)(135),lamdaOut => P(2)(391));
U_G3392: entity G port map(lamdaA => P(3)(264),lamdaB => P(3)(392),s => s(3)(136),lamdaOut => P(2)(392));
U_G3393: entity G port map(lamdaA => P(3)(265),lamdaB => P(3)(393),s => s(3)(137),lamdaOut => P(2)(393));
U_G3394: entity G port map(lamdaA => P(3)(266),lamdaB => P(3)(394),s => s(3)(138),lamdaOut => P(2)(394));
U_G3395: entity G port map(lamdaA => P(3)(267),lamdaB => P(3)(395),s => s(3)(139),lamdaOut => P(2)(395));
U_G3396: entity G port map(lamdaA => P(3)(268),lamdaB => P(3)(396),s => s(3)(140),lamdaOut => P(2)(396));
U_G3397: entity G port map(lamdaA => P(3)(269),lamdaB => P(3)(397),s => s(3)(141),lamdaOut => P(2)(397));
U_G3398: entity G port map(lamdaA => P(3)(270),lamdaB => P(3)(398),s => s(3)(142),lamdaOut => P(2)(398));
U_G3399: entity G port map(lamdaA => P(3)(271),lamdaB => P(3)(399),s => s(3)(143),lamdaOut => P(2)(399));
U_G3400: entity G port map(lamdaA => P(3)(272),lamdaB => P(3)(400),s => s(3)(144),lamdaOut => P(2)(400));
U_G3401: entity G port map(lamdaA => P(3)(273),lamdaB => P(3)(401),s => s(3)(145),lamdaOut => P(2)(401));
U_G3402: entity G port map(lamdaA => P(3)(274),lamdaB => P(3)(402),s => s(3)(146),lamdaOut => P(2)(402));
U_G3403: entity G port map(lamdaA => P(3)(275),lamdaB => P(3)(403),s => s(3)(147),lamdaOut => P(2)(403));
U_G3404: entity G port map(lamdaA => P(3)(276),lamdaB => P(3)(404),s => s(3)(148),lamdaOut => P(2)(404));
U_G3405: entity G port map(lamdaA => P(3)(277),lamdaB => P(3)(405),s => s(3)(149),lamdaOut => P(2)(405));
U_G3406: entity G port map(lamdaA => P(3)(278),lamdaB => P(3)(406),s => s(3)(150),lamdaOut => P(2)(406));
U_G3407: entity G port map(lamdaA => P(3)(279),lamdaB => P(3)(407),s => s(3)(151),lamdaOut => P(2)(407));
U_G3408: entity G port map(lamdaA => P(3)(280),lamdaB => P(3)(408),s => s(3)(152),lamdaOut => P(2)(408));
U_G3409: entity G port map(lamdaA => P(3)(281),lamdaB => P(3)(409),s => s(3)(153),lamdaOut => P(2)(409));
U_G3410: entity G port map(lamdaA => P(3)(282),lamdaB => P(3)(410),s => s(3)(154),lamdaOut => P(2)(410));
U_G3411: entity G port map(lamdaA => P(3)(283),lamdaB => P(3)(411),s => s(3)(155),lamdaOut => P(2)(411));
U_G3412: entity G port map(lamdaA => P(3)(284),lamdaB => P(3)(412),s => s(3)(156),lamdaOut => P(2)(412));
U_G3413: entity G port map(lamdaA => P(3)(285),lamdaB => P(3)(413),s => s(3)(157),lamdaOut => P(2)(413));
U_G3414: entity G port map(lamdaA => P(3)(286),lamdaB => P(3)(414),s => s(3)(158),lamdaOut => P(2)(414));
U_G3415: entity G port map(lamdaA => P(3)(287),lamdaB => P(3)(415),s => s(3)(159),lamdaOut => P(2)(415));
U_G3416: entity G port map(lamdaA => P(3)(288),lamdaB => P(3)(416),s => s(3)(160),lamdaOut => P(2)(416));
U_G3417: entity G port map(lamdaA => P(3)(289),lamdaB => P(3)(417),s => s(3)(161),lamdaOut => P(2)(417));
U_G3418: entity G port map(lamdaA => P(3)(290),lamdaB => P(3)(418),s => s(3)(162),lamdaOut => P(2)(418));
U_G3419: entity G port map(lamdaA => P(3)(291),lamdaB => P(3)(419),s => s(3)(163),lamdaOut => P(2)(419));
U_G3420: entity G port map(lamdaA => P(3)(292),lamdaB => P(3)(420),s => s(3)(164),lamdaOut => P(2)(420));
U_G3421: entity G port map(lamdaA => P(3)(293),lamdaB => P(3)(421),s => s(3)(165),lamdaOut => P(2)(421));
U_G3422: entity G port map(lamdaA => P(3)(294),lamdaB => P(3)(422),s => s(3)(166),lamdaOut => P(2)(422));
U_G3423: entity G port map(lamdaA => P(3)(295),lamdaB => P(3)(423),s => s(3)(167),lamdaOut => P(2)(423));
U_G3424: entity G port map(lamdaA => P(3)(296),lamdaB => P(3)(424),s => s(3)(168),lamdaOut => P(2)(424));
U_G3425: entity G port map(lamdaA => P(3)(297),lamdaB => P(3)(425),s => s(3)(169),lamdaOut => P(2)(425));
U_G3426: entity G port map(lamdaA => P(3)(298),lamdaB => P(3)(426),s => s(3)(170),lamdaOut => P(2)(426));
U_G3427: entity G port map(lamdaA => P(3)(299),lamdaB => P(3)(427),s => s(3)(171),lamdaOut => P(2)(427));
U_G3428: entity G port map(lamdaA => P(3)(300),lamdaB => P(3)(428),s => s(3)(172),lamdaOut => P(2)(428));
U_G3429: entity G port map(lamdaA => P(3)(301),lamdaB => P(3)(429),s => s(3)(173),lamdaOut => P(2)(429));
U_G3430: entity G port map(lamdaA => P(3)(302),lamdaB => P(3)(430),s => s(3)(174),lamdaOut => P(2)(430));
U_G3431: entity G port map(lamdaA => P(3)(303),lamdaB => P(3)(431),s => s(3)(175),lamdaOut => P(2)(431));
U_G3432: entity G port map(lamdaA => P(3)(304),lamdaB => P(3)(432),s => s(3)(176),lamdaOut => P(2)(432));
U_G3433: entity G port map(lamdaA => P(3)(305),lamdaB => P(3)(433),s => s(3)(177),lamdaOut => P(2)(433));
U_G3434: entity G port map(lamdaA => P(3)(306),lamdaB => P(3)(434),s => s(3)(178),lamdaOut => P(2)(434));
U_G3435: entity G port map(lamdaA => P(3)(307),lamdaB => P(3)(435),s => s(3)(179),lamdaOut => P(2)(435));
U_G3436: entity G port map(lamdaA => P(3)(308),lamdaB => P(3)(436),s => s(3)(180),lamdaOut => P(2)(436));
U_G3437: entity G port map(lamdaA => P(3)(309),lamdaB => P(3)(437),s => s(3)(181),lamdaOut => P(2)(437));
U_G3438: entity G port map(lamdaA => P(3)(310),lamdaB => P(3)(438),s => s(3)(182),lamdaOut => P(2)(438));
U_G3439: entity G port map(lamdaA => P(3)(311),lamdaB => P(3)(439),s => s(3)(183),lamdaOut => P(2)(439));
U_G3440: entity G port map(lamdaA => P(3)(312),lamdaB => P(3)(440),s => s(3)(184),lamdaOut => P(2)(440));
U_G3441: entity G port map(lamdaA => P(3)(313),lamdaB => P(3)(441),s => s(3)(185),lamdaOut => P(2)(441));
U_G3442: entity G port map(lamdaA => P(3)(314),lamdaB => P(3)(442),s => s(3)(186),lamdaOut => P(2)(442));
U_G3443: entity G port map(lamdaA => P(3)(315),lamdaB => P(3)(443),s => s(3)(187),lamdaOut => P(2)(443));
U_G3444: entity G port map(lamdaA => P(3)(316),lamdaB => P(3)(444),s => s(3)(188),lamdaOut => P(2)(444));
U_G3445: entity G port map(lamdaA => P(3)(317),lamdaB => P(3)(445),s => s(3)(189),lamdaOut => P(2)(445));
U_G3446: entity G port map(lamdaA => P(3)(318),lamdaB => P(3)(446),s => s(3)(190),lamdaOut => P(2)(446));
U_G3447: entity G port map(lamdaA => P(3)(319),lamdaB => P(3)(447),s => s(3)(191),lamdaOut => P(2)(447));
U_G3448: entity G port map(lamdaA => P(3)(320),lamdaB => P(3)(448),s => s(3)(192),lamdaOut => P(2)(448));
U_G3449: entity G port map(lamdaA => P(3)(321),lamdaB => P(3)(449),s => s(3)(193),lamdaOut => P(2)(449));
U_G3450: entity G port map(lamdaA => P(3)(322),lamdaB => P(3)(450),s => s(3)(194),lamdaOut => P(2)(450));
U_G3451: entity G port map(lamdaA => P(3)(323),lamdaB => P(3)(451),s => s(3)(195),lamdaOut => P(2)(451));
U_G3452: entity G port map(lamdaA => P(3)(324),lamdaB => P(3)(452),s => s(3)(196),lamdaOut => P(2)(452));
U_G3453: entity G port map(lamdaA => P(3)(325),lamdaB => P(3)(453),s => s(3)(197),lamdaOut => P(2)(453));
U_G3454: entity G port map(lamdaA => P(3)(326),lamdaB => P(3)(454),s => s(3)(198),lamdaOut => P(2)(454));
U_G3455: entity G port map(lamdaA => P(3)(327),lamdaB => P(3)(455),s => s(3)(199),lamdaOut => P(2)(455));
U_G3456: entity G port map(lamdaA => P(3)(328),lamdaB => P(3)(456),s => s(3)(200),lamdaOut => P(2)(456));
U_G3457: entity G port map(lamdaA => P(3)(329),lamdaB => P(3)(457),s => s(3)(201),lamdaOut => P(2)(457));
U_G3458: entity G port map(lamdaA => P(3)(330),lamdaB => P(3)(458),s => s(3)(202),lamdaOut => P(2)(458));
U_G3459: entity G port map(lamdaA => P(3)(331),lamdaB => P(3)(459),s => s(3)(203),lamdaOut => P(2)(459));
U_G3460: entity G port map(lamdaA => P(3)(332),lamdaB => P(3)(460),s => s(3)(204),lamdaOut => P(2)(460));
U_G3461: entity G port map(lamdaA => P(3)(333),lamdaB => P(3)(461),s => s(3)(205),lamdaOut => P(2)(461));
U_G3462: entity G port map(lamdaA => P(3)(334),lamdaB => P(3)(462),s => s(3)(206),lamdaOut => P(2)(462));
U_G3463: entity G port map(lamdaA => P(3)(335),lamdaB => P(3)(463),s => s(3)(207),lamdaOut => P(2)(463));
U_G3464: entity G port map(lamdaA => P(3)(336),lamdaB => P(3)(464),s => s(3)(208),lamdaOut => P(2)(464));
U_G3465: entity G port map(lamdaA => P(3)(337),lamdaB => P(3)(465),s => s(3)(209),lamdaOut => P(2)(465));
U_G3466: entity G port map(lamdaA => P(3)(338),lamdaB => P(3)(466),s => s(3)(210),lamdaOut => P(2)(466));
U_G3467: entity G port map(lamdaA => P(3)(339),lamdaB => P(3)(467),s => s(3)(211),lamdaOut => P(2)(467));
U_G3468: entity G port map(lamdaA => P(3)(340),lamdaB => P(3)(468),s => s(3)(212),lamdaOut => P(2)(468));
U_G3469: entity G port map(lamdaA => P(3)(341),lamdaB => P(3)(469),s => s(3)(213),lamdaOut => P(2)(469));
U_G3470: entity G port map(lamdaA => P(3)(342),lamdaB => P(3)(470),s => s(3)(214),lamdaOut => P(2)(470));
U_G3471: entity G port map(lamdaA => P(3)(343),lamdaB => P(3)(471),s => s(3)(215),lamdaOut => P(2)(471));
U_G3472: entity G port map(lamdaA => P(3)(344),lamdaB => P(3)(472),s => s(3)(216),lamdaOut => P(2)(472));
U_G3473: entity G port map(lamdaA => P(3)(345),lamdaB => P(3)(473),s => s(3)(217),lamdaOut => P(2)(473));
U_G3474: entity G port map(lamdaA => P(3)(346),lamdaB => P(3)(474),s => s(3)(218),lamdaOut => P(2)(474));
U_G3475: entity G port map(lamdaA => P(3)(347),lamdaB => P(3)(475),s => s(3)(219),lamdaOut => P(2)(475));
U_G3476: entity G port map(lamdaA => P(3)(348),lamdaB => P(3)(476),s => s(3)(220),lamdaOut => P(2)(476));
U_G3477: entity G port map(lamdaA => P(3)(349),lamdaB => P(3)(477),s => s(3)(221),lamdaOut => P(2)(477));
U_G3478: entity G port map(lamdaA => P(3)(350),lamdaB => P(3)(478),s => s(3)(222),lamdaOut => P(2)(478));
U_G3479: entity G port map(lamdaA => P(3)(351),lamdaB => P(3)(479),s => s(3)(223),lamdaOut => P(2)(479));
U_G3480: entity G port map(lamdaA => P(3)(352),lamdaB => P(3)(480),s => s(3)(224),lamdaOut => P(2)(480));
U_G3481: entity G port map(lamdaA => P(3)(353),lamdaB => P(3)(481),s => s(3)(225),lamdaOut => P(2)(481));
U_G3482: entity G port map(lamdaA => P(3)(354),lamdaB => P(3)(482),s => s(3)(226),lamdaOut => P(2)(482));
U_G3483: entity G port map(lamdaA => P(3)(355),lamdaB => P(3)(483),s => s(3)(227),lamdaOut => P(2)(483));
U_G3484: entity G port map(lamdaA => P(3)(356),lamdaB => P(3)(484),s => s(3)(228),lamdaOut => P(2)(484));
U_G3485: entity G port map(lamdaA => P(3)(357),lamdaB => P(3)(485),s => s(3)(229),lamdaOut => P(2)(485));
U_G3486: entity G port map(lamdaA => P(3)(358),lamdaB => P(3)(486),s => s(3)(230),lamdaOut => P(2)(486));
U_G3487: entity G port map(lamdaA => P(3)(359),lamdaB => P(3)(487),s => s(3)(231),lamdaOut => P(2)(487));
U_G3488: entity G port map(lamdaA => P(3)(360),lamdaB => P(3)(488),s => s(3)(232),lamdaOut => P(2)(488));
U_G3489: entity G port map(lamdaA => P(3)(361),lamdaB => P(3)(489),s => s(3)(233),lamdaOut => P(2)(489));
U_G3490: entity G port map(lamdaA => P(3)(362),lamdaB => P(3)(490),s => s(3)(234),lamdaOut => P(2)(490));
U_G3491: entity G port map(lamdaA => P(3)(363),lamdaB => P(3)(491),s => s(3)(235),lamdaOut => P(2)(491));
U_G3492: entity G port map(lamdaA => P(3)(364),lamdaB => P(3)(492),s => s(3)(236),lamdaOut => P(2)(492));
U_G3493: entity G port map(lamdaA => P(3)(365),lamdaB => P(3)(493),s => s(3)(237),lamdaOut => P(2)(493));
U_G3494: entity G port map(lamdaA => P(3)(366),lamdaB => P(3)(494),s => s(3)(238),lamdaOut => P(2)(494));
U_G3495: entity G port map(lamdaA => P(3)(367),lamdaB => P(3)(495),s => s(3)(239),lamdaOut => P(2)(495));
U_G3496: entity G port map(lamdaA => P(3)(368),lamdaB => P(3)(496),s => s(3)(240),lamdaOut => P(2)(496));
U_G3497: entity G port map(lamdaA => P(3)(369),lamdaB => P(3)(497),s => s(3)(241),lamdaOut => P(2)(497));
U_G3498: entity G port map(lamdaA => P(3)(370),lamdaB => P(3)(498),s => s(3)(242),lamdaOut => P(2)(498));
U_G3499: entity G port map(lamdaA => P(3)(371),lamdaB => P(3)(499),s => s(3)(243),lamdaOut => P(2)(499));
U_G3500: entity G port map(lamdaA => P(3)(372),lamdaB => P(3)(500),s => s(3)(244),lamdaOut => P(2)(500));
U_G3501: entity G port map(lamdaA => P(3)(373),lamdaB => P(3)(501),s => s(3)(245),lamdaOut => P(2)(501));
U_G3502: entity G port map(lamdaA => P(3)(374),lamdaB => P(3)(502),s => s(3)(246),lamdaOut => P(2)(502));
U_G3503: entity G port map(lamdaA => P(3)(375),lamdaB => P(3)(503),s => s(3)(247),lamdaOut => P(2)(503));
U_G3504: entity G port map(lamdaA => P(3)(376),lamdaB => P(3)(504),s => s(3)(248),lamdaOut => P(2)(504));
U_G3505: entity G port map(lamdaA => P(3)(377),lamdaB => P(3)(505),s => s(3)(249),lamdaOut => P(2)(505));
U_G3506: entity G port map(lamdaA => P(3)(378),lamdaB => P(3)(506),s => s(3)(250),lamdaOut => P(2)(506));
U_G3507: entity G port map(lamdaA => P(3)(379),lamdaB => P(3)(507),s => s(3)(251),lamdaOut => P(2)(507));
U_G3508: entity G port map(lamdaA => P(3)(380),lamdaB => P(3)(508),s => s(3)(252),lamdaOut => P(2)(508));
U_G3509: entity G port map(lamdaA => P(3)(381),lamdaB => P(3)(509),s => s(3)(253),lamdaOut => P(2)(509));
U_G3510: entity G port map(lamdaA => P(3)(382),lamdaB => P(3)(510),s => s(3)(254),lamdaOut => P(2)(510));
U_G3511: entity G port map(lamdaA => P(3)(383),lamdaB => P(3)(511),s => s(3)(255),lamdaOut => P(2)(511));
U_F3512: entity F port map(lamdaA => P(3)(512),lamdaB => P(3)(640),lamdaOut => P(2)(512));
U_F3513: entity F port map(lamdaA => P(3)(513),lamdaB => P(3)(641),lamdaOut => P(2)(513));
U_F3514: entity F port map(lamdaA => P(3)(514),lamdaB => P(3)(642),lamdaOut => P(2)(514));
U_F3515: entity F port map(lamdaA => P(3)(515),lamdaB => P(3)(643),lamdaOut => P(2)(515));
U_F3516: entity F port map(lamdaA => P(3)(516),lamdaB => P(3)(644),lamdaOut => P(2)(516));
U_F3517: entity F port map(lamdaA => P(3)(517),lamdaB => P(3)(645),lamdaOut => P(2)(517));
U_F3518: entity F port map(lamdaA => P(3)(518),lamdaB => P(3)(646),lamdaOut => P(2)(518));
U_F3519: entity F port map(lamdaA => P(3)(519),lamdaB => P(3)(647),lamdaOut => P(2)(519));
U_F3520: entity F port map(lamdaA => P(3)(520),lamdaB => P(3)(648),lamdaOut => P(2)(520));
U_F3521: entity F port map(lamdaA => P(3)(521),lamdaB => P(3)(649),lamdaOut => P(2)(521));
U_F3522: entity F port map(lamdaA => P(3)(522),lamdaB => P(3)(650),lamdaOut => P(2)(522));
U_F3523: entity F port map(lamdaA => P(3)(523),lamdaB => P(3)(651),lamdaOut => P(2)(523));
U_F3524: entity F port map(lamdaA => P(3)(524),lamdaB => P(3)(652),lamdaOut => P(2)(524));
U_F3525: entity F port map(lamdaA => P(3)(525),lamdaB => P(3)(653),lamdaOut => P(2)(525));
U_F3526: entity F port map(lamdaA => P(3)(526),lamdaB => P(3)(654),lamdaOut => P(2)(526));
U_F3527: entity F port map(lamdaA => P(3)(527),lamdaB => P(3)(655),lamdaOut => P(2)(527));
U_F3528: entity F port map(lamdaA => P(3)(528),lamdaB => P(3)(656),lamdaOut => P(2)(528));
U_F3529: entity F port map(lamdaA => P(3)(529),lamdaB => P(3)(657),lamdaOut => P(2)(529));
U_F3530: entity F port map(lamdaA => P(3)(530),lamdaB => P(3)(658),lamdaOut => P(2)(530));
U_F3531: entity F port map(lamdaA => P(3)(531),lamdaB => P(3)(659),lamdaOut => P(2)(531));
U_F3532: entity F port map(lamdaA => P(3)(532),lamdaB => P(3)(660),lamdaOut => P(2)(532));
U_F3533: entity F port map(lamdaA => P(3)(533),lamdaB => P(3)(661),lamdaOut => P(2)(533));
U_F3534: entity F port map(lamdaA => P(3)(534),lamdaB => P(3)(662),lamdaOut => P(2)(534));
U_F3535: entity F port map(lamdaA => P(3)(535),lamdaB => P(3)(663),lamdaOut => P(2)(535));
U_F3536: entity F port map(lamdaA => P(3)(536),lamdaB => P(3)(664),lamdaOut => P(2)(536));
U_F3537: entity F port map(lamdaA => P(3)(537),lamdaB => P(3)(665),lamdaOut => P(2)(537));
U_F3538: entity F port map(lamdaA => P(3)(538),lamdaB => P(3)(666),lamdaOut => P(2)(538));
U_F3539: entity F port map(lamdaA => P(3)(539),lamdaB => P(3)(667),lamdaOut => P(2)(539));
U_F3540: entity F port map(lamdaA => P(3)(540),lamdaB => P(3)(668),lamdaOut => P(2)(540));
U_F3541: entity F port map(lamdaA => P(3)(541),lamdaB => P(3)(669),lamdaOut => P(2)(541));
U_F3542: entity F port map(lamdaA => P(3)(542),lamdaB => P(3)(670),lamdaOut => P(2)(542));
U_F3543: entity F port map(lamdaA => P(3)(543),lamdaB => P(3)(671),lamdaOut => P(2)(543));
U_F3544: entity F port map(lamdaA => P(3)(544),lamdaB => P(3)(672),lamdaOut => P(2)(544));
U_F3545: entity F port map(lamdaA => P(3)(545),lamdaB => P(3)(673),lamdaOut => P(2)(545));
U_F3546: entity F port map(lamdaA => P(3)(546),lamdaB => P(3)(674),lamdaOut => P(2)(546));
U_F3547: entity F port map(lamdaA => P(3)(547),lamdaB => P(3)(675),lamdaOut => P(2)(547));
U_F3548: entity F port map(lamdaA => P(3)(548),lamdaB => P(3)(676),lamdaOut => P(2)(548));
U_F3549: entity F port map(lamdaA => P(3)(549),lamdaB => P(3)(677),lamdaOut => P(2)(549));
U_F3550: entity F port map(lamdaA => P(3)(550),lamdaB => P(3)(678),lamdaOut => P(2)(550));
U_F3551: entity F port map(lamdaA => P(3)(551),lamdaB => P(3)(679),lamdaOut => P(2)(551));
U_F3552: entity F port map(lamdaA => P(3)(552),lamdaB => P(3)(680),lamdaOut => P(2)(552));
U_F3553: entity F port map(lamdaA => P(3)(553),lamdaB => P(3)(681),lamdaOut => P(2)(553));
U_F3554: entity F port map(lamdaA => P(3)(554),lamdaB => P(3)(682),lamdaOut => P(2)(554));
U_F3555: entity F port map(lamdaA => P(3)(555),lamdaB => P(3)(683),lamdaOut => P(2)(555));
U_F3556: entity F port map(lamdaA => P(3)(556),lamdaB => P(3)(684),lamdaOut => P(2)(556));
U_F3557: entity F port map(lamdaA => P(3)(557),lamdaB => P(3)(685),lamdaOut => P(2)(557));
U_F3558: entity F port map(lamdaA => P(3)(558),lamdaB => P(3)(686),lamdaOut => P(2)(558));
U_F3559: entity F port map(lamdaA => P(3)(559),lamdaB => P(3)(687),lamdaOut => P(2)(559));
U_F3560: entity F port map(lamdaA => P(3)(560),lamdaB => P(3)(688),lamdaOut => P(2)(560));
U_F3561: entity F port map(lamdaA => P(3)(561),lamdaB => P(3)(689),lamdaOut => P(2)(561));
U_F3562: entity F port map(lamdaA => P(3)(562),lamdaB => P(3)(690),lamdaOut => P(2)(562));
U_F3563: entity F port map(lamdaA => P(3)(563),lamdaB => P(3)(691),lamdaOut => P(2)(563));
U_F3564: entity F port map(lamdaA => P(3)(564),lamdaB => P(3)(692),lamdaOut => P(2)(564));
U_F3565: entity F port map(lamdaA => P(3)(565),lamdaB => P(3)(693),lamdaOut => P(2)(565));
U_F3566: entity F port map(lamdaA => P(3)(566),lamdaB => P(3)(694),lamdaOut => P(2)(566));
U_F3567: entity F port map(lamdaA => P(3)(567),lamdaB => P(3)(695),lamdaOut => P(2)(567));
U_F3568: entity F port map(lamdaA => P(3)(568),lamdaB => P(3)(696),lamdaOut => P(2)(568));
U_F3569: entity F port map(lamdaA => P(3)(569),lamdaB => P(3)(697),lamdaOut => P(2)(569));
U_F3570: entity F port map(lamdaA => P(3)(570),lamdaB => P(3)(698),lamdaOut => P(2)(570));
U_F3571: entity F port map(lamdaA => P(3)(571),lamdaB => P(3)(699),lamdaOut => P(2)(571));
U_F3572: entity F port map(lamdaA => P(3)(572),lamdaB => P(3)(700),lamdaOut => P(2)(572));
U_F3573: entity F port map(lamdaA => P(3)(573),lamdaB => P(3)(701),lamdaOut => P(2)(573));
U_F3574: entity F port map(lamdaA => P(3)(574),lamdaB => P(3)(702),lamdaOut => P(2)(574));
U_F3575: entity F port map(lamdaA => P(3)(575),lamdaB => P(3)(703),lamdaOut => P(2)(575));
U_F3576: entity F port map(lamdaA => P(3)(576),lamdaB => P(3)(704),lamdaOut => P(2)(576));
U_F3577: entity F port map(lamdaA => P(3)(577),lamdaB => P(3)(705),lamdaOut => P(2)(577));
U_F3578: entity F port map(lamdaA => P(3)(578),lamdaB => P(3)(706),lamdaOut => P(2)(578));
U_F3579: entity F port map(lamdaA => P(3)(579),lamdaB => P(3)(707),lamdaOut => P(2)(579));
U_F3580: entity F port map(lamdaA => P(3)(580),lamdaB => P(3)(708),lamdaOut => P(2)(580));
U_F3581: entity F port map(lamdaA => P(3)(581),lamdaB => P(3)(709),lamdaOut => P(2)(581));
U_F3582: entity F port map(lamdaA => P(3)(582),lamdaB => P(3)(710),lamdaOut => P(2)(582));
U_F3583: entity F port map(lamdaA => P(3)(583),lamdaB => P(3)(711),lamdaOut => P(2)(583));
U_F3584: entity F port map(lamdaA => P(3)(584),lamdaB => P(3)(712),lamdaOut => P(2)(584));
U_F3585: entity F port map(lamdaA => P(3)(585),lamdaB => P(3)(713),lamdaOut => P(2)(585));
U_F3586: entity F port map(lamdaA => P(3)(586),lamdaB => P(3)(714),lamdaOut => P(2)(586));
U_F3587: entity F port map(lamdaA => P(3)(587),lamdaB => P(3)(715),lamdaOut => P(2)(587));
U_F3588: entity F port map(lamdaA => P(3)(588),lamdaB => P(3)(716),lamdaOut => P(2)(588));
U_F3589: entity F port map(lamdaA => P(3)(589),lamdaB => P(3)(717),lamdaOut => P(2)(589));
U_F3590: entity F port map(lamdaA => P(3)(590),lamdaB => P(3)(718),lamdaOut => P(2)(590));
U_F3591: entity F port map(lamdaA => P(3)(591),lamdaB => P(3)(719),lamdaOut => P(2)(591));
U_F3592: entity F port map(lamdaA => P(3)(592),lamdaB => P(3)(720),lamdaOut => P(2)(592));
U_F3593: entity F port map(lamdaA => P(3)(593),lamdaB => P(3)(721),lamdaOut => P(2)(593));
U_F3594: entity F port map(lamdaA => P(3)(594),lamdaB => P(3)(722),lamdaOut => P(2)(594));
U_F3595: entity F port map(lamdaA => P(3)(595),lamdaB => P(3)(723),lamdaOut => P(2)(595));
U_F3596: entity F port map(lamdaA => P(3)(596),lamdaB => P(3)(724),lamdaOut => P(2)(596));
U_F3597: entity F port map(lamdaA => P(3)(597),lamdaB => P(3)(725),lamdaOut => P(2)(597));
U_F3598: entity F port map(lamdaA => P(3)(598),lamdaB => P(3)(726),lamdaOut => P(2)(598));
U_F3599: entity F port map(lamdaA => P(3)(599),lamdaB => P(3)(727),lamdaOut => P(2)(599));
U_F3600: entity F port map(lamdaA => P(3)(600),lamdaB => P(3)(728),lamdaOut => P(2)(600));
U_F3601: entity F port map(lamdaA => P(3)(601),lamdaB => P(3)(729),lamdaOut => P(2)(601));
U_F3602: entity F port map(lamdaA => P(3)(602),lamdaB => P(3)(730),lamdaOut => P(2)(602));
U_F3603: entity F port map(lamdaA => P(3)(603),lamdaB => P(3)(731),lamdaOut => P(2)(603));
U_F3604: entity F port map(lamdaA => P(3)(604),lamdaB => P(3)(732),lamdaOut => P(2)(604));
U_F3605: entity F port map(lamdaA => P(3)(605),lamdaB => P(3)(733),lamdaOut => P(2)(605));
U_F3606: entity F port map(lamdaA => P(3)(606),lamdaB => P(3)(734),lamdaOut => P(2)(606));
U_F3607: entity F port map(lamdaA => P(3)(607),lamdaB => P(3)(735),lamdaOut => P(2)(607));
U_F3608: entity F port map(lamdaA => P(3)(608),lamdaB => P(3)(736),lamdaOut => P(2)(608));
U_F3609: entity F port map(lamdaA => P(3)(609),lamdaB => P(3)(737),lamdaOut => P(2)(609));
U_F3610: entity F port map(lamdaA => P(3)(610),lamdaB => P(3)(738),lamdaOut => P(2)(610));
U_F3611: entity F port map(lamdaA => P(3)(611),lamdaB => P(3)(739),lamdaOut => P(2)(611));
U_F3612: entity F port map(lamdaA => P(3)(612),lamdaB => P(3)(740),lamdaOut => P(2)(612));
U_F3613: entity F port map(lamdaA => P(3)(613),lamdaB => P(3)(741),lamdaOut => P(2)(613));
U_F3614: entity F port map(lamdaA => P(3)(614),lamdaB => P(3)(742),lamdaOut => P(2)(614));
U_F3615: entity F port map(lamdaA => P(3)(615),lamdaB => P(3)(743),lamdaOut => P(2)(615));
U_F3616: entity F port map(lamdaA => P(3)(616),lamdaB => P(3)(744),lamdaOut => P(2)(616));
U_F3617: entity F port map(lamdaA => P(3)(617),lamdaB => P(3)(745),lamdaOut => P(2)(617));
U_F3618: entity F port map(lamdaA => P(3)(618),lamdaB => P(3)(746),lamdaOut => P(2)(618));
U_F3619: entity F port map(lamdaA => P(3)(619),lamdaB => P(3)(747),lamdaOut => P(2)(619));
U_F3620: entity F port map(lamdaA => P(3)(620),lamdaB => P(3)(748),lamdaOut => P(2)(620));
U_F3621: entity F port map(lamdaA => P(3)(621),lamdaB => P(3)(749),lamdaOut => P(2)(621));
U_F3622: entity F port map(lamdaA => P(3)(622),lamdaB => P(3)(750),lamdaOut => P(2)(622));
U_F3623: entity F port map(lamdaA => P(3)(623),lamdaB => P(3)(751),lamdaOut => P(2)(623));
U_F3624: entity F port map(lamdaA => P(3)(624),lamdaB => P(3)(752),lamdaOut => P(2)(624));
U_F3625: entity F port map(lamdaA => P(3)(625),lamdaB => P(3)(753),lamdaOut => P(2)(625));
U_F3626: entity F port map(lamdaA => P(3)(626),lamdaB => P(3)(754),lamdaOut => P(2)(626));
U_F3627: entity F port map(lamdaA => P(3)(627),lamdaB => P(3)(755),lamdaOut => P(2)(627));
U_F3628: entity F port map(lamdaA => P(3)(628),lamdaB => P(3)(756),lamdaOut => P(2)(628));
U_F3629: entity F port map(lamdaA => P(3)(629),lamdaB => P(3)(757),lamdaOut => P(2)(629));
U_F3630: entity F port map(lamdaA => P(3)(630),lamdaB => P(3)(758),lamdaOut => P(2)(630));
U_F3631: entity F port map(lamdaA => P(3)(631),lamdaB => P(3)(759),lamdaOut => P(2)(631));
U_F3632: entity F port map(lamdaA => P(3)(632),lamdaB => P(3)(760),lamdaOut => P(2)(632));
U_F3633: entity F port map(lamdaA => P(3)(633),lamdaB => P(3)(761),lamdaOut => P(2)(633));
U_F3634: entity F port map(lamdaA => P(3)(634),lamdaB => P(3)(762),lamdaOut => P(2)(634));
U_F3635: entity F port map(lamdaA => P(3)(635),lamdaB => P(3)(763),lamdaOut => P(2)(635));
U_F3636: entity F port map(lamdaA => P(3)(636),lamdaB => P(3)(764),lamdaOut => P(2)(636));
U_F3637: entity F port map(lamdaA => P(3)(637),lamdaB => P(3)(765),lamdaOut => P(2)(637));
U_F3638: entity F port map(lamdaA => P(3)(638),lamdaB => P(3)(766),lamdaOut => P(2)(638));
U_F3639: entity F port map(lamdaA => P(3)(639),lamdaB => P(3)(767),lamdaOut => P(2)(639));
U_G3640: entity G port map(lamdaA => P(3)(512),lamdaB => P(3)(640),s => s(3)(256),lamdaOut => P(2)(640));
U_G3641: entity G port map(lamdaA => P(3)(513),lamdaB => P(3)(641),s => s(3)(257),lamdaOut => P(2)(641));
U_G3642: entity G port map(lamdaA => P(3)(514),lamdaB => P(3)(642),s => s(3)(258),lamdaOut => P(2)(642));
U_G3643: entity G port map(lamdaA => P(3)(515),lamdaB => P(3)(643),s => s(3)(259),lamdaOut => P(2)(643));
U_G3644: entity G port map(lamdaA => P(3)(516),lamdaB => P(3)(644),s => s(3)(260),lamdaOut => P(2)(644));
U_G3645: entity G port map(lamdaA => P(3)(517),lamdaB => P(3)(645),s => s(3)(261),lamdaOut => P(2)(645));
U_G3646: entity G port map(lamdaA => P(3)(518),lamdaB => P(3)(646),s => s(3)(262),lamdaOut => P(2)(646));
U_G3647: entity G port map(lamdaA => P(3)(519),lamdaB => P(3)(647),s => s(3)(263),lamdaOut => P(2)(647));
U_G3648: entity G port map(lamdaA => P(3)(520),lamdaB => P(3)(648),s => s(3)(264),lamdaOut => P(2)(648));
U_G3649: entity G port map(lamdaA => P(3)(521),lamdaB => P(3)(649),s => s(3)(265),lamdaOut => P(2)(649));
U_G3650: entity G port map(lamdaA => P(3)(522),lamdaB => P(3)(650),s => s(3)(266),lamdaOut => P(2)(650));
U_G3651: entity G port map(lamdaA => P(3)(523),lamdaB => P(3)(651),s => s(3)(267),lamdaOut => P(2)(651));
U_G3652: entity G port map(lamdaA => P(3)(524),lamdaB => P(3)(652),s => s(3)(268),lamdaOut => P(2)(652));
U_G3653: entity G port map(lamdaA => P(3)(525),lamdaB => P(3)(653),s => s(3)(269),lamdaOut => P(2)(653));
U_G3654: entity G port map(lamdaA => P(3)(526),lamdaB => P(3)(654),s => s(3)(270),lamdaOut => P(2)(654));
U_G3655: entity G port map(lamdaA => P(3)(527),lamdaB => P(3)(655),s => s(3)(271),lamdaOut => P(2)(655));
U_G3656: entity G port map(lamdaA => P(3)(528),lamdaB => P(3)(656),s => s(3)(272),lamdaOut => P(2)(656));
U_G3657: entity G port map(lamdaA => P(3)(529),lamdaB => P(3)(657),s => s(3)(273),lamdaOut => P(2)(657));
U_G3658: entity G port map(lamdaA => P(3)(530),lamdaB => P(3)(658),s => s(3)(274),lamdaOut => P(2)(658));
U_G3659: entity G port map(lamdaA => P(3)(531),lamdaB => P(3)(659),s => s(3)(275),lamdaOut => P(2)(659));
U_G3660: entity G port map(lamdaA => P(3)(532),lamdaB => P(3)(660),s => s(3)(276),lamdaOut => P(2)(660));
U_G3661: entity G port map(lamdaA => P(3)(533),lamdaB => P(3)(661),s => s(3)(277),lamdaOut => P(2)(661));
U_G3662: entity G port map(lamdaA => P(3)(534),lamdaB => P(3)(662),s => s(3)(278),lamdaOut => P(2)(662));
U_G3663: entity G port map(lamdaA => P(3)(535),lamdaB => P(3)(663),s => s(3)(279),lamdaOut => P(2)(663));
U_G3664: entity G port map(lamdaA => P(3)(536),lamdaB => P(3)(664),s => s(3)(280),lamdaOut => P(2)(664));
U_G3665: entity G port map(lamdaA => P(3)(537),lamdaB => P(3)(665),s => s(3)(281),lamdaOut => P(2)(665));
U_G3666: entity G port map(lamdaA => P(3)(538),lamdaB => P(3)(666),s => s(3)(282),lamdaOut => P(2)(666));
U_G3667: entity G port map(lamdaA => P(3)(539),lamdaB => P(3)(667),s => s(3)(283),lamdaOut => P(2)(667));
U_G3668: entity G port map(lamdaA => P(3)(540),lamdaB => P(3)(668),s => s(3)(284),lamdaOut => P(2)(668));
U_G3669: entity G port map(lamdaA => P(3)(541),lamdaB => P(3)(669),s => s(3)(285),lamdaOut => P(2)(669));
U_G3670: entity G port map(lamdaA => P(3)(542),lamdaB => P(3)(670),s => s(3)(286),lamdaOut => P(2)(670));
U_G3671: entity G port map(lamdaA => P(3)(543),lamdaB => P(3)(671),s => s(3)(287),lamdaOut => P(2)(671));
U_G3672: entity G port map(lamdaA => P(3)(544),lamdaB => P(3)(672),s => s(3)(288),lamdaOut => P(2)(672));
U_G3673: entity G port map(lamdaA => P(3)(545),lamdaB => P(3)(673),s => s(3)(289),lamdaOut => P(2)(673));
U_G3674: entity G port map(lamdaA => P(3)(546),lamdaB => P(3)(674),s => s(3)(290),lamdaOut => P(2)(674));
U_G3675: entity G port map(lamdaA => P(3)(547),lamdaB => P(3)(675),s => s(3)(291),lamdaOut => P(2)(675));
U_G3676: entity G port map(lamdaA => P(3)(548),lamdaB => P(3)(676),s => s(3)(292),lamdaOut => P(2)(676));
U_G3677: entity G port map(lamdaA => P(3)(549),lamdaB => P(3)(677),s => s(3)(293),lamdaOut => P(2)(677));
U_G3678: entity G port map(lamdaA => P(3)(550),lamdaB => P(3)(678),s => s(3)(294),lamdaOut => P(2)(678));
U_G3679: entity G port map(lamdaA => P(3)(551),lamdaB => P(3)(679),s => s(3)(295),lamdaOut => P(2)(679));
U_G3680: entity G port map(lamdaA => P(3)(552),lamdaB => P(3)(680),s => s(3)(296),lamdaOut => P(2)(680));
U_G3681: entity G port map(lamdaA => P(3)(553),lamdaB => P(3)(681),s => s(3)(297),lamdaOut => P(2)(681));
U_G3682: entity G port map(lamdaA => P(3)(554),lamdaB => P(3)(682),s => s(3)(298),lamdaOut => P(2)(682));
U_G3683: entity G port map(lamdaA => P(3)(555),lamdaB => P(3)(683),s => s(3)(299),lamdaOut => P(2)(683));
U_G3684: entity G port map(lamdaA => P(3)(556),lamdaB => P(3)(684),s => s(3)(300),lamdaOut => P(2)(684));
U_G3685: entity G port map(lamdaA => P(3)(557),lamdaB => P(3)(685),s => s(3)(301),lamdaOut => P(2)(685));
U_G3686: entity G port map(lamdaA => P(3)(558),lamdaB => P(3)(686),s => s(3)(302),lamdaOut => P(2)(686));
U_G3687: entity G port map(lamdaA => P(3)(559),lamdaB => P(3)(687),s => s(3)(303),lamdaOut => P(2)(687));
U_G3688: entity G port map(lamdaA => P(3)(560),lamdaB => P(3)(688),s => s(3)(304),lamdaOut => P(2)(688));
U_G3689: entity G port map(lamdaA => P(3)(561),lamdaB => P(3)(689),s => s(3)(305),lamdaOut => P(2)(689));
U_G3690: entity G port map(lamdaA => P(3)(562),lamdaB => P(3)(690),s => s(3)(306),lamdaOut => P(2)(690));
U_G3691: entity G port map(lamdaA => P(3)(563),lamdaB => P(3)(691),s => s(3)(307),lamdaOut => P(2)(691));
U_G3692: entity G port map(lamdaA => P(3)(564),lamdaB => P(3)(692),s => s(3)(308),lamdaOut => P(2)(692));
U_G3693: entity G port map(lamdaA => P(3)(565),lamdaB => P(3)(693),s => s(3)(309),lamdaOut => P(2)(693));
U_G3694: entity G port map(lamdaA => P(3)(566),lamdaB => P(3)(694),s => s(3)(310),lamdaOut => P(2)(694));
U_G3695: entity G port map(lamdaA => P(3)(567),lamdaB => P(3)(695),s => s(3)(311),lamdaOut => P(2)(695));
U_G3696: entity G port map(lamdaA => P(3)(568),lamdaB => P(3)(696),s => s(3)(312),lamdaOut => P(2)(696));
U_G3697: entity G port map(lamdaA => P(3)(569),lamdaB => P(3)(697),s => s(3)(313),lamdaOut => P(2)(697));
U_G3698: entity G port map(lamdaA => P(3)(570),lamdaB => P(3)(698),s => s(3)(314),lamdaOut => P(2)(698));
U_G3699: entity G port map(lamdaA => P(3)(571),lamdaB => P(3)(699),s => s(3)(315),lamdaOut => P(2)(699));
U_G3700: entity G port map(lamdaA => P(3)(572),lamdaB => P(3)(700),s => s(3)(316),lamdaOut => P(2)(700));
U_G3701: entity G port map(lamdaA => P(3)(573),lamdaB => P(3)(701),s => s(3)(317),lamdaOut => P(2)(701));
U_G3702: entity G port map(lamdaA => P(3)(574),lamdaB => P(3)(702),s => s(3)(318),lamdaOut => P(2)(702));
U_G3703: entity G port map(lamdaA => P(3)(575),lamdaB => P(3)(703),s => s(3)(319),lamdaOut => P(2)(703));
U_G3704: entity G port map(lamdaA => P(3)(576),lamdaB => P(3)(704),s => s(3)(320),lamdaOut => P(2)(704));
U_G3705: entity G port map(lamdaA => P(3)(577),lamdaB => P(3)(705),s => s(3)(321),lamdaOut => P(2)(705));
U_G3706: entity G port map(lamdaA => P(3)(578),lamdaB => P(3)(706),s => s(3)(322),lamdaOut => P(2)(706));
U_G3707: entity G port map(lamdaA => P(3)(579),lamdaB => P(3)(707),s => s(3)(323),lamdaOut => P(2)(707));
U_G3708: entity G port map(lamdaA => P(3)(580),lamdaB => P(3)(708),s => s(3)(324),lamdaOut => P(2)(708));
U_G3709: entity G port map(lamdaA => P(3)(581),lamdaB => P(3)(709),s => s(3)(325),lamdaOut => P(2)(709));
U_G3710: entity G port map(lamdaA => P(3)(582),lamdaB => P(3)(710),s => s(3)(326),lamdaOut => P(2)(710));
U_G3711: entity G port map(lamdaA => P(3)(583),lamdaB => P(3)(711),s => s(3)(327),lamdaOut => P(2)(711));
U_G3712: entity G port map(lamdaA => P(3)(584),lamdaB => P(3)(712),s => s(3)(328),lamdaOut => P(2)(712));
U_G3713: entity G port map(lamdaA => P(3)(585),lamdaB => P(3)(713),s => s(3)(329),lamdaOut => P(2)(713));
U_G3714: entity G port map(lamdaA => P(3)(586),lamdaB => P(3)(714),s => s(3)(330),lamdaOut => P(2)(714));
U_G3715: entity G port map(lamdaA => P(3)(587),lamdaB => P(3)(715),s => s(3)(331),lamdaOut => P(2)(715));
U_G3716: entity G port map(lamdaA => P(3)(588),lamdaB => P(3)(716),s => s(3)(332),lamdaOut => P(2)(716));
U_G3717: entity G port map(lamdaA => P(3)(589),lamdaB => P(3)(717),s => s(3)(333),lamdaOut => P(2)(717));
U_G3718: entity G port map(lamdaA => P(3)(590),lamdaB => P(3)(718),s => s(3)(334),lamdaOut => P(2)(718));
U_G3719: entity G port map(lamdaA => P(3)(591),lamdaB => P(3)(719),s => s(3)(335),lamdaOut => P(2)(719));
U_G3720: entity G port map(lamdaA => P(3)(592),lamdaB => P(3)(720),s => s(3)(336),lamdaOut => P(2)(720));
U_G3721: entity G port map(lamdaA => P(3)(593),lamdaB => P(3)(721),s => s(3)(337),lamdaOut => P(2)(721));
U_G3722: entity G port map(lamdaA => P(3)(594),lamdaB => P(3)(722),s => s(3)(338),lamdaOut => P(2)(722));
U_G3723: entity G port map(lamdaA => P(3)(595),lamdaB => P(3)(723),s => s(3)(339),lamdaOut => P(2)(723));
U_G3724: entity G port map(lamdaA => P(3)(596),lamdaB => P(3)(724),s => s(3)(340),lamdaOut => P(2)(724));
U_G3725: entity G port map(lamdaA => P(3)(597),lamdaB => P(3)(725),s => s(3)(341),lamdaOut => P(2)(725));
U_G3726: entity G port map(lamdaA => P(3)(598),lamdaB => P(3)(726),s => s(3)(342),lamdaOut => P(2)(726));
U_G3727: entity G port map(lamdaA => P(3)(599),lamdaB => P(3)(727),s => s(3)(343),lamdaOut => P(2)(727));
U_G3728: entity G port map(lamdaA => P(3)(600),lamdaB => P(3)(728),s => s(3)(344),lamdaOut => P(2)(728));
U_G3729: entity G port map(lamdaA => P(3)(601),lamdaB => P(3)(729),s => s(3)(345),lamdaOut => P(2)(729));
U_G3730: entity G port map(lamdaA => P(3)(602),lamdaB => P(3)(730),s => s(3)(346),lamdaOut => P(2)(730));
U_G3731: entity G port map(lamdaA => P(3)(603),lamdaB => P(3)(731),s => s(3)(347),lamdaOut => P(2)(731));
U_G3732: entity G port map(lamdaA => P(3)(604),lamdaB => P(3)(732),s => s(3)(348),lamdaOut => P(2)(732));
U_G3733: entity G port map(lamdaA => P(3)(605),lamdaB => P(3)(733),s => s(3)(349),lamdaOut => P(2)(733));
U_G3734: entity G port map(lamdaA => P(3)(606),lamdaB => P(3)(734),s => s(3)(350),lamdaOut => P(2)(734));
U_G3735: entity G port map(lamdaA => P(3)(607),lamdaB => P(3)(735),s => s(3)(351),lamdaOut => P(2)(735));
U_G3736: entity G port map(lamdaA => P(3)(608),lamdaB => P(3)(736),s => s(3)(352),lamdaOut => P(2)(736));
U_G3737: entity G port map(lamdaA => P(3)(609),lamdaB => P(3)(737),s => s(3)(353),lamdaOut => P(2)(737));
U_G3738: entity G port map(lamdaA => P(3)(610),lamdaB => P(3)(738),s => s(3)(354),lamdaOut => P(2)(738));
U_G3739: entity G port map(lamdaA => P(3)(611),lamdaB => P(3)(739),s => s(3)(355),lamdaOut => P(2)(739));
U_G3740: entity G port map(lamdaA => P(3)(612),lamdaB => P(3)(740),s => s(3)(356),lamdaOut => P(2)(740));
U_G3741: entity G port map(lamdaA => P(3)(613),lamdaB => P(3)(741),s => s(3)(357),lamdaOut => P(2)(741));
U_G3742: entity G port map(lamdaA => P(3)(614),lamdaB => P(3)(742),s => s(3)(358),lamdaOut => P(2)(742));
U_G3743: entity G port map(lamdaA => P(3)(615),lamdaB => P(3)(743),s => s(3)(359),lamdaOut => P(2)(743));
U_G3744: entity G port map(lamdaA => P(3)(616),lamdaB => P(3)(744),s => s(3)(360),lamdaOut => P(2)(744));
U_G3745: entity G port map(lamdaA => P(3)(617),lamdaB => P(3)(745),s => s(3)(361),lamdaOut => P(2)(745));
U_G3746: entity G port map(lamdaA => P(3)(618),lamdaB => P(3)(746),s => s(3)(362),lamdaOut => P(2)(746));
U_G3747: entity G port map(lamdaA => P(3)(619),lamdaB => P(3)(747),s => s(3)(363),lamdaOut => P(2)(747));
U_G3748: entity G port map(lamdaA => P(3)(620),lamdaB => P(3)(748),s => s(3)(364),lamdaOut => P(2)(748));
U_G3749: entity G port map(lamdaA => P(3)(621),lamdaB => P(3)(749),s => s(3)(365),lamdaOut => P(2)(749));
U_G3750: entity G port map(lamdaA => P(3)(622),lamdaB => P(3)(750),s => s(3)(366),lamdaOut => P(2)(750));
U_G3751: entity G port map(lamdaA => P(3)(623),lamdaB => P(3)(751),s => s(3)(367),lamdaOut => P(2)(751));
U_G3752: entity G port map(lamdaA => P(3)(624),lamdaB => P(3)(752),s => s(3)(368),lamdaOut => P(2)(752));
U_G3753: entity G port map(lamdaA => P(3)(625),lamdaB => P(3)(753),s => s(3)(369),lamdaOut => P(2)(753));
U_G3754: entity G port map(lamdaA => P(3)(626),lamdaB => P(3)(754),s => s(3)(370),lamdaOut => P(2)(754));
U_G3755: entity G port map(lamdaA => P(3)(627),lamdaB => P(3)(755),s => s(3)(371),lamdaOut => P(2)(755));
U_G3756: entity G port map(lamdaA => P(3)(628),lamdaB => P(3)(756),s => s(3)(372),lamdaOut => P(2)(756));
U_G3757: entity G port map(lamdaA => P(3)(629),lamdaB => P(3)(757),s => s(3)(373),lamdaOut => P(2)(757));
U_G3758: entity G port map(lamdaA => P(3)(630),lamdaB => P(3)(758),s => s(3)(374),lamdaOut => P(2)(758));
U_G3759: entity G port map(lamdaA => P(3)(631),lamdaB => P(3)(759),s => s(3)(375),lamdaOut => P(2)(759));
U_G3760: entity G port map(lamdaA => P(3)(632),lamdaB => P(3)(760),s => s(3)(376),lamdaOut => P(2)(760));
U_G3761: entity G port map(lamdaA => P(3)(633),lamdaB => P(3)(761),s => s(3)(377),lamdaOut => P(2)(761));
U_G3762: entity G port map(lamdaA => P(3)(634),lamdaB => P(3)(762),s => s(3)(378),lamdaOut => P(2)(762));
U_G3763: entity G port map(lamdaA => P(3)(635),lamdaB => P(3)(763),s => s(3)(379),lamdaOut => P(2)(763));
U_G3764: entity G port map(lamdaA => P(3)(636),lamdaB => P(3)(764),s => s(3)(380),lamdaOut => P(2)(764));
U_G3765: entity G port map(lamdaA => P(3)(637),lamdaB => P(3)(765),s => s(3)(381),lamdaOut => P(2)(765));
U_G3766: entity G port map(lamdaA => P(3)(638),lamdaB => P(3)(766),s => s(3)(382),lamdaOut => P(2)(766));
U_G3767: entity G port map(lamdaA => P(3)(639),lamdaB => P(3)(767),s => s(3)(383),lamdaOut => P(2)(767));
U_F3768: entity F port map(lamdaA => P(3)(768),lamdaB => P(3)(896),lamdaOut => P(2)(768));
U_F3769: entity F port map(lamdaA => P(3)(769),lamdaB => P(3)(897),lamdaOut => P(2)(769));
U_F3770: entity F port map(lamdaA => P(3)(770),lamdaB => P(3)(898),lamdaOut => P(2)(770));
U_F3771: entity F port map(lamdaA => P(3)(771),lamdaB => P(3)(899),lamdaOut => P(2)(771));
U_F3772: entity F port map(lamdaA => P(3)(772),lamdaB => P(3)(900),lamdaOut => P(2)(772));
U_F3773: entity F port map(lamdaA => P(3)(773),lamdaB => P(3)(901),lamdaOut => P(2)(773));
U_F3774: entity F port map(lamdaA => P(3)(774),lamdaB => P(3)(902),lamdaOut => P(2)(774));
U_F3775: entity F port map(lamdaA => P(3)(775),lamdaB => P(3)(903),lamdaOut => P(2)(775));
U_F3776: entity F port map(lamdaA => P(3)(776),lamdaB => P(3)(904),lamdaOut => P(2)(776));
U_F3777: entity F port map(lamdaA => P(3)(777),lamdaB => P(3)(905),lamdaOut => P(2)(777));
U_F3778: entity F port map(lamdaA => P(3)(778),lamdaB => P(3)(906),lamdaOut => P(2)(778));
U_F3779: entity F port map(lamdaA => P(3)(779),lamdaB => P(3)(907),lamdaOut => P(2)(779));
U_F3780: entity F port map(lamdaA => P(3)(780),lamdaB => P(3)(908),lamdaOut => P(2)(780));
U_F3781: entity F port map(lamdaA => P(3)(781),lamdaB => P(3)(909),lamdaOut => P(2)(781));
U_F3782: entity F port map(lamdaA => P(3)(782),lamdaB => P(3)(910),lamdaOut => P(2)(782));
U_F3783: entity F port map(lamdaA => P(3)(783),lamdaB => P(3)(911),lamdaOut => P(2)(783));
U_F3784: entity F port map(lamdaA => P(3)(784),lamdaB => P(3)(912),lamdaOut => P(2)(784));
U_F3785: entity F port map(lamdaA => P(3)(785),lamdaB => P(3)(913),lamdaOut => P(2)(785));
U_F3786: entity F port map(lamdaA => P(3)(786),lamdaB => P(3)(914),lamdaOut => P(2)(786));
U_F3787: entity F port map(lamdaA => P(3)(787),lamdaB => P(3)(915),lamdaOut => P(2)(787));
U_F3788: entity F port map(lamdaA => P(3)(788),lamdaB => P(3)(916),lamdaOut => P(2)(788));
U_F3789: entity F port map(lamdaA => P(3)(789),lamdaB => P(3)(917),lamdaOut => P(2)(789));
U_F3790: entity F port map(lamdaA => P(3)(790),lamdaB => P(3)(918),lamdaOut => P(2)(790));
U_F3791: entity F port map(lamdaA => P(3)(791),lamdaB => P(3)(919),lamdaOut => P(2)(791));
U_F3792: entity F port map(lamdaA => P(3)(792),lamdaB => P(3)(920),lamdaOut => P(2)(792));
U_F3793: entity F port map(lamdaA => P(3)(793),lamdaB => P(3)(921),lamdaOut => P(2)(793));
U_F3794: entity F port map(lamdaA => P(3)(794),lamdaB => P(3)(922),lamdaOut => P(2)(794));
U_F3795: entity F port map(lamdaA => P(3)(795),lamdaB => P(3)(923),lamdaOut => P(2)(795));
U_F3796: entity F port map(lamdaA => P(3)(796),lamdaB => P(3)(924),lamdaOut => P(2)(796));
U_F3797: entity F port map(lamdaA => P(3)(797),lamdaB => P(3)(925),lamdaOut => P(2)(797));
U_F3798: entity F port map(lamdaA => P(3)(798),lamdaB => P(3)(926),lamdaOut => P(2)(798));
U_F3799: entity F port map(lamdaA => P(3)(799),lamdaB => P(3)(927),lamdaOut => P(2)(799));
U_F3800: entity F port map(lamdaA => P(3)(800),lamdaB => P(3)(928),lamdaOut => P(2)(800));
U_F3801: entity F port map(lamdaA => P(3)(801),lamdaB => P(3)(929),lamdaOut => P(2)(801));
U_F3802: entity F port map(lamdaA => P(3)(802),lamdaB => P(3)(930),lamdaOut => P(2)(802));
U_F3803: entity F port map(lamdaA => P(3)(803),lamdaB => P(3)(931),lamdaOut => P(2)(803));
U_F3804: entity F port map(lamdaA => P(3)(804),lamdaB => P(3)(932),lamdaOut => P(2)(804));
U_F3805: entity F port map(lamdaA => P(3)(805),lamdaB => P(3)(933),lamdaOut => P(2)(805));
U_F3806: entity F port map(lamdaA => P(3)(806),lamdaB => P(3)(934),lamdaOut => P(2)(806));
U_F3807: entity F port map(lamdaA => P(3)(807),lamdaB => P(3)(935),lamdaOut => P(2)(807));
U_F3808: entity F port map(lamdaA => P(3)(808),lamdaB => P(3)(936),lamdaOut => P(2)(808));
U_F3809: entity F port map(lamdaA => P(3)(809),lamdaB => P(3)(937),lamdaOut => P(2)(809));
U_F3810: entity F port map(lamdaA => P(3)(810),lamdaB => P(3)(938),lamdaOut => P(2)(810));
U_F3811: entity F port map(lamdaA => P(3)(811),lamdaB => P(3)(939),lamdaOut => P(2)(811));
U_F3812: entity F port map(lamdaA => P(3)(812),lamdaB => P(3)(940),lamdaOut => P(2)(812));
U_F3813: entity F port map(lamdaA => P(3)(813),lamdaB => P(3)(941),lamdaOut => P(2)(813));
U_F3814: entity F port map(lamdaA => P(3)(814),lamdaB => P(3)(942),lamdaOut => P(2)(814));
U_F3815: entity F port map(lamdaA => P(3)(815),lamdaB => P(3)(943),lamdaOut => P(2)(815));
U_F3816: entity F port map(lamdaA => P(3)(816),lamdaB => P(3)(944),lamdaOut => P(2)(816));
U_F3817: entity F port map(lamdaA => P(3)(817),lamdaB => P(3)(945),lamdaOut => P(2)(817));
U_F3818: entity F port map(lamdaA => P(3)(818),lamdaB => P(3)(946),lamdaOut => P(2)(818));
U_F3819: entity F port map(lamdaA => P(3)(819),lamdaB => P(3)(947),lamdaOut => P(2)(819));
U_F3820: entity F port map(lamdaA => P(3)(820),lamdaB => P(3)(948),lamdaOut => P(2)(820));
U_F3821: entity F port map(lamdaA => P(3)(821),lamdaB => P(3)(949),lamdaOut => P(2)(821));
U_F3822: entity F port map(lamdaA => P(3)(822),lamdaB => P(3)(950),lamdaOut => P(2)(822));
U_F3823: entity F port map(lamdaA => P(3)(823),lamdaB => P(3)(951),lamdaOut => P(2)(823));
U_F3824: entity F port map(lamdaA => P(3)(824),lamdaB => P(3)(952),lamdaOut => P(2)(824));
U_F3825: entity F port map(lamdaA => P(3)(825),lamdaB => P(3)(953),lamdaOut => P(2)(825));
U_F3826: entity F port map(lamdaA => P(3)(826),lamdaB => P(3)(954),lamdaOut => P(2)(826));
U_F3827: entity F port map(lamdaA => P(3)(827),lamdaB => P(3)(955),lamdaOut => P(2)(827));
U_F3828: entity F port map(lamdaA => P(3)(828),lamdaB => P(3)(956),lamdaOut => P(2)(828));
U_F3829: entity F port map(lamdaA => P(3)(829),lamdaB => P(3)(957),lamdaOut => P(2)(829));
U_F3830: entity F port map(lamdaA => P(3)(830),lamdaB => P(3)(958),lamdaOut => P(2)(830));
U_F3831: entity F port map(lamdaA => P(3)(831),lamdaB => P(3)(959),lamdaOut => P(2)(831));
U_F3832: entity F port map(lamdaA => P(3)(832),lamdaB => P(3)(960),lamdaOut => P(2)(832));
U_F3833: entity F port map(lamdaA => P(3)(833),lamdaB => P(3)(961),lamdaOut => P(2)(833));
U_F3834: entity F port map(lamdaA => P(3)(834),lamdaB => P(3)(962),lamdaOut => P(2)(834));
U_F3835: entity F port map(lamdaA => P(3)(835),lamdaB => P(3)(963),lamdaOut => P(2)(835));
U_F3836: entity F port map(lamdaA => P(3)(836),lamdaB => P(3)(964),lamdaOut => P(2)(836));
U_F3837: entity F port map(lamdaA => P(3)(837),lamdaB => P(3)(965),lamdaOut => P(2)(837));
U_F3838: entity F port map(lamdaA => P(3)(838),lamdaB => P(3)(966),lamdaOut => P(2)(838));
U_F3839: entity F port map(lamdaA => P(3)(839),lamdaB => P(3)(967),lamdaOut => P(2)(839));
U_F3840: entity F port map(lamdaA => P(3)(840),lamdaB => P(3)(968),lamdaOut => P(2)(840));
U_F3841: entity F port map(lamdaA => P(3)(841),lamdaB => P(3)(969),lamdaOut => P(2)(841));
U_F3842: entity F port map(lamdaA => P(3)(842),lamdaB => P(3)(970),lamdaOut => P(2)(842));
U_F3843: entity F port map(lamdaA => P(3)(843),lamdaB => P(3)(971),lamdaOut => P(2)(843));
U_F3844: entity F port map(lamdaA => P(3)(844),lamdaB => P(3)(972),lamdaOut => P(2)(844));
U_F3845: entity F port map(lamdaA => P(3)(845),lamdaB => P(3)(973),lamdaOut => P(2)(845));
U_F3846: entity F port map(lamdaA => P(3)(846),lamdaB => P(3)(974),lamdaOut => P(2)(846));
U_F3847: entity F port map(lamdaA => P(3)(847),lamdaB => P(3)(975),lamdaOut => P(2)(847));
U_F3848: entity F port map(lamdaA => P(3)(848),lamdaB => P(3)(976),lamdaOut => P(2)(848));
U_F3849: entity F port map(lamdaA => P(3)(849),lamdaB => P(3)(977),lamdaOut => P(2)(849));
U_F3850: entity F port map(lamdaA => P(3)(850),lamdaB => P(3)(978),lamdaOut => P(2)(850));
U_F3851: entity F port map(lamdaA => P(3)(851),lamdaB => P(3)(979),lamdaOut => P(2)(851));
U_F3852: entity F port map(lamdaA => P(3)(852),lamdaB => P(3)(980),lamdaOut => P(2)(852));
U_F3853: entity F port map(lamdaA => P(3)(853),lamdaB => P(3)(981),lamdaOut => P(2)(853));
U_F3854: entity F port map(lamdaA => P(3)(854),lamdaB => P(3)(982),lamdaOut => P(2)(854));
U_F3855: entity F port map(lamdaA => P(3)(855),lamdaB => P(3)(983),lamdaOut => P(2)(855));
U_F3856: entity F port map(lamdaA => P(3)(856),lamdaB => P(3)(984),lamdaOut => P(2)(856));
U_F3857: entity F port map(lamdaA => P(3)(857),lamdaB => P(3)(985),lamdaOut => P(2)(857));
U_F3858: entity F port map(lamdaA => P(3)(858),lamdaB => P(3)(986),lamdaOut => P(2)(858));
U_F3859: entity F port map(lamdaA => P(3)(859),lamdaB => P(3)(987),lamdaOut => P(2)(859));
U_F3860: entity F port map(lamdaA => P(3)(860),lamdaB => P(3)(988),lamdaOut => P(2)(860));
U_F3861: entity F port map(lamdaA => P(3)(861),lamdaB => P(3)(989),lamdaOut => P(2)(861));
U_F3862: entity F port map(lamdaA => P(3)(862),lamdaB => P(3)(990),lamdaOut => P(2)(862));
U_F3863: entity F port map(lamdaA => P(3)(863),lamdaB => P(3)(991),lamdaOut => P(2)(863));
U_F3864: entity F port map(lamdaA => P(3)(864),lamdaB => P(3)(992),lamdaOut => P(2)(864));
U_F3865: entity F port map(lamdaA => P(3)(865),lamdaB => P(3)(993),lamdaOut => P(2)(865));
U_F3866: entity F port map(lamdaA => P(3)(866),lamdaB => P(3)(994),lamdaOut => P(2)(866));
U_F3867: entity F port map(lamdaA => P(3)(867),lamdaB => P(3)(995),lamdaOut => P(2)(867));
U_F3868: entity F port map(lamdaA => P(3)(868),lamdaB => P(3)(996),lamdaOut => P(2)(868));
U_F3869: entity F port map(lamdaA => P(3)(869),lamdaB => P(3)(997),lamdaOut => P(2)(869));
U_F3870: entity F port map(lamdaA => P(3)(870),lamdaB => P(3)(998),lamdaOut => P(2)(870));
U_F3871: entity F port map(lamdaA => P(3)(871),lamdaB => P(3)(999),lamdaOut => P(2)(871));
U_F3872: entity F port map(lamdaA => P(3)(872),lamdaB => P(3)(1000),lamdaOut => P(2)(872));
U_F3873: entity F port map(lamdaA => P(3)(873),lamdaB => P(3)(1001),lamdaOut => P(2)(873));
U_F3874: entity F port map(lamdaA => P(3)(874),lamdaB => P(3)(1002),lamdaOut => P(2)(874));
U_F3875: entity F port map(lamdaA => P(3)(875),lamdaB => P(3)(1003),lamdaOut => P(2)(875));
U_F3876: entity F port map(lamdaA => P(3)(876),lamdaB => P(3)(1004),lamdaOut => P(2)(876));
U_F3877: entity F port map(lamdaA => P(3)(877),lamdaB => P(3)(1005),lamdaOut => P(2)(877));
U_F3878: entity F port map(lamdaA => P(3)(878),lamdaB => P(3)(1006),lamdaOut => P(2)(878));
U_F3879: entity F port map(lamdaA => P(3)(879),lamdaB => P(3)(1007),lamdaOut => P(2)(879));
U_F3880: entity F port map(lamdaA => P(3)(880),lamdaB => P(3)(1008),lamdaOut => P(2)(880));
U_F3881: entity F port map(lamdaA => P(3)(881),lamdaB => P(3)(1009),lamdaOut => P(2)(881));
U_F3882: entity F port map(lamdaA => P(3)(882),lamdaB => P(3)(1010),lamdaOut => P(2)(882));
U_F3883: entity F port map(lamdaA => P(3)(883),lamdaB => P(3)(1011),lamdaOut => P(2)(883));
U_F3884: entity F port map(lamdaA => P(3)(884),lamdaB => P(3)(1012),lamdaOut => P(2)(884));
U_F3885: entity F port map(lamdaA => P(3)(885),lamdaB => P(3)(1013),lamdaOut => P(2)(885));
U_F3886: entity F port map(lamdaA => P(3)(886),lamdaB => P(3)(1014),lamdaOut => P(2)(886));
U_F3887: entity F port map(lamdaA => P(3)(887),lamdaB => P(3)(1015),lamdaOut => P(2)(887));
U_F3888: entity F port map(lamdaA => P(3)(888),lamdaB => P(3)(1016),lamdaOut => P(2)(888));
U_F3889: entity F port map(lamdaA => P(3)(889),lamdaB => P(3)(1017),lamdaOut => P(2)(889));
U_F3890: entity F port map(lamdaA => P(3)(890),lamdaB => P(3)(1018),lamdaOut => P(2)(890));
U_F3891: entity F port map(lamdaA => P(3)(891),lamdaB => P(3)(1019),lamdaOut => P(2)(891));
U_F3892: entity F port map(lamdaA => P(3)(892),lamdaB => P(3)(1020),lamdaOut => P(2)(892));
U_F3893: entity F port map(lamdaA => P(3)(893),lamdaB => P(3)(1021),lamdaOut => P(2)(893));
U_F3894: entity F port map(lamdaA => P(3)(894),lamdaB => P(3)(1022),lamdaOut => P(2)(894));
U_F3895: entity F port map(lamdaA => P(3)(895),lamdaB => P(3)(1023),lamdaOut => P(2)(895));
U_G3896: entity G port map(lamdaA => P(3)(768),lamdaB => P(3)(896),s => s(3)(384),lamdaOut => P(2)(896));
U_G3897: entity G port map(lamdaA => P(3)(769),lamdaB => P(3)(897),s => s(3)(385),lamdaOut => P(2)(897));
U_G3898: entity G port map(lamdaA => P(3)(770),lamdaB => P(3)(898),s => s(3)(386),lamdaOut => P(2)(898));
U_G3899: entity G port map(lamdaA => P(3)(771),lamdaB => P(3)(899),s => s(3)(387),lamdaOut => P(2)(899));
U_G3900: entity G port map(lamdaA => P(3)(772),lamdaB => P(3)(900),s => s(3)(388),lamdaOut => P(2)(900));
U_G3901: entity G port map(lamdaA => P(3)(773),lamdaB => P(3)(901),s => s(3)(389),lamdaOut => P(2)(901));
U_G3902: entity G port map(lamdaA => P(3)(774),lamdaB => P(3)(902),s => s(3)(390),lamdaOut => P(2)(902));
U_G3903: entity G port map(lamdaA => P(3)(775),lamdaB => P(3)(903),s => s(3)(391),lamdaOut => P(2)(903));
U_G3904: entity G port map(lamdaA => P(3)(776),lamdaB => P(3)(904),s => s(3)(392),lamdaOut => P(2)(904));
U_G3905: entity G port map(lamdaA => P(3)(777),lamdaB => P(3)(905),s => s(3)(393),lamdaOut => P(2)(905));
U_G3906: entity G port map(lamdaA => P(3)(778),lamdaB => P(3)(906),s => s(3)(394),lamdaOut => P(2)(906));
U_G3907: entity G port map(lamdaA => P(3)(779),lamdaB => P(3)(907),s => s(3)(395),lamdaOut => P(2)(907));
U_G3908: entity G port map(lamdaA => P(3)(780),lamdaB => P(3)(908),s => s(3)(396),lamdaOut => P(2)(908));
U_G3909: entity G port map(lamdaA => P(3)(781),lamdaB => P(3)(909),s => s(3)(397),lamdaOut => P(2)(909));
U_G3910: entity G port map(lamdaA => P(3)(782),lamdaB => P(3)(910),s => s(3)(398),lamdaOut => P(2)(910));
U_G3911: entity G port map(lamdaA => P(3)(783),lamdaB => P(3)(911),s => s(3)(399),lamdaOut => P(2)(911));
U_G3912: entity G port map(lamdaA => P(3)(784),lamdaB => P(3)(912),s => s(3)(400),lamdaOut => P(2)(912));
U_G3913: entity G port map(lamdaA => P(3)(785),lamdaB => P(3)(913),s => s(3)(401),lamdaOut => P(2)(913));
U_G3914: entity G port map(lamdaA => P(3)(786),lamdaB => P(3)(914),s => s(3)(402),lamdaOut => P(2)(914));
U_G3915: entity G port map(lamdaA => P(3)(787),lamdaB => P(3)(915),s => s(3)(403),lamdaOut => P(2)(915));
U_G3916: entity G port map(lamdaA => P(3)(788),lamdaB => P(3)(916),s => s(3)(404),lamdaOut => P(2)(916));
U_G3917: entity G port map(lamdaA => P(3)(789),lamdaB => P(3)(917),s => s(3)(405),lamdaOut => P(2)(917));
U_G3918: entity G port map(lamdaA => P(3)(790),lamdaB => P(3)(918),s => s(3)(406),lamdaOut => P(2)(918));
U_G3919: entity G port map(lamdaA => P(3)(791),lamdaB => P(3)(919),s => s(3)(407),lamdaOut => P(2)(919));
U_G3920: entity G port map(lamdaA => P(3)(792),lamdaB => P(3)(920),s => s(3)(408),lamdaOut => P(2)(920));
U_G3921: entity G port map(lamdaA => P(3)(793),lamdaB => P(3)(921),s => s(3)(409),lamdaOut => P(2)(921));
U_G3922: entity G port map(lamdaA => P(3)(794),lamdaB => P(3)(922),s => s(3)(410),lamdaOut => P(2)(922));
U_G3923: entity G port map(lamdaA => P(3)(795),lamdaB => P(3)(923),s => s(3)(411),lamdaOut => P(2)(923));
U_G3924: entity G port map(lamdaA => P(3)(796),lamdaB => P(3)(924),s => s(3)(412),lamdaOut => P(2)(924));
U_G3925: entity G port map(lamdaA => P(3)(797),lamdaB => P(3)(925),s => s(3)(413),lamdaOut => P(2)(925));
U_G3926: entity G port map(lamdaA => P(3)(798),lamdaB => P(3)(926),s => s(3)(414),lamdaOut => P(2)(926));
U_G3927: entity G port map(lamdaA => P(3)(799),lamdaB => P(3)(927),s => s(3)(415),lamdaOut => P(2)(927));
U_G3928: entity G port map(lamdaA => P(3)(800),lamdaB => P(3)(928),s => s(3)(416),lamdaOut => P(2)(928));
U_G3929: entity G port map(lamdaA => P(3)(801),lamdaB => P(3)(929),s => s(3)(417),lamdaOut => P(2)(929));
U_G3930: entity G port map(lamdaA => P(3)(802),lamdaB => P(3)(930),s => s(3)(418),lamdaOut => P(2)(930));
U_G3931: entity G port map(lamdaA => P(3)(803),lamdaB => P(3)(931),s => s(3)(419),lamdaOut => P(2)(931));
U_G3932: entity G port map(lamdaA => P(3)(804),lamdaB => P(3)(932),s => s(3)(420),lamdaOut => P(2)(932));
U_G3933: entity G port map(lamdaA => P(3)(805),lamdaB => P(3)(933),s => s(3)(421),lamdaOut => P(2)(933));
U_G3934: entity G port map(lamdaA => P(3)(806),lamdaB => P(3)(934),s => s(3)(422),lamdaOut => P(2)(934));
U_G3935: entity G port map(lamdaA => P(3)(807),lamdaB => P(3)(935),s => s(3)(423),lamdaOut => P(2)(935));
U_G3936: entity G port map(lamdaA => P(3)(808),lamdaB => P(3)(936),s => s(3)(424),lamdaOut => P(2)(936));
U_G3937: entity G port map(lamdaA => P(3)(809),lamdaB => P(3)(937),s => s(3)(425),lamdaOut => P(2)(937));
U_G3938: entity G port map(lamdaA => P(3)(810),lamdaB => P(3)(938),s => s(3)(426),lamdaOut => P(2)(938));
U_G3939: entity G port map(lamdaA => P(3)(811),lamdaB => P(3)(939),s => s(3)(427),lamdaOut => P(2)(939));
U_G3940: entity G port map(lamdaA => P(3)(812),lamdaB => P(3)(940),s => s(3)(428),lamdaOut => P(2)(940));
U_G3941: entity G port map(lamdaA => P(3)(813),lamdaB => P(3)(941),s => s(3)(429),lamdaOut => P(2)(941));
U_G3942: entity G port map(lamdaA => P(3)(814),lamdaB => P(3)(942),s => s(3)(430),lamdaOut => P(2)(942));
U_G3943: entity G port map(lamdaA => P(3)(815),lamdaB => P(3)(943),s => s(3)(431),lamdaOut => P(2)(943));
U_G3944: entity G port map(lamdaA => P(3)(816),lamdaB => P(3)(944),s => s(3)(432),lamdaOut => P(2)(944));
U_G3945: entity G port map(lamdaA => P(3)(817),lamdaB => P(3)(945),s => s(3)(433),lamdaOut => P(2)(945));
U_G3946: entity G port map(lamdaA => P(3)(818),lamdaB => P(3)(946),s => s(3)(434),lamdaOut => P(2)(946));
U_G3947: entity G port map(lamdaA => P(3)(819),lamdaB => P(3)(947),s => s(3)(435),lamdaOut => P(2)(947));
U_G3948: entity G port map(lamdaA => P(3)(820),lamdaB => P(3)(948),s => s(3)(436),lamdaOut => P(2)(948));
U_G3949: entity G port map(lamdaA => P(3)(821),lamdaB => P(3)(949),s => s(3)(437),lamdaOut => P(2)(949));
U_G3950: entity G port map(lamdaA => P(3)(822),lamdaB => P(3)(950),s => s(3)(438),lamdaOut => P(2)(950));
U_G3951: entity G port map(lamdaA => P(3)(823),lamdaB => P(3)(951),s => s(3)(439),lamdaOut => P(2)(951));
U_G3952: entity G port map(lamdaA => P(3)(824),lamdaB => P(3)(952),s => s(3)(440),lamdaOut => P(2)(952));
U_G3953: entity G port map(lamdaA => P(3)(825),lamdaB => P(3)(953),s => s(3)(441),lamdaOut => P(2)(953));
U_G3954: entity G port map(lamdaA => P(3)(826),lamdaB => P(3)(954),s => s(3)(442),lamdaOut => P(2)(954));
U_G3955: entity G port map(lamdaA => P(3)(827),lamdaB => P(3)(955),s => s(3)(443),lamdaOut => P(2)(955));
U_G3956: entity G port map(lamdaA => P(3)(828),lamdaB => P(3)(956),s => s(3)(444),lamdaOut => P(2)(956));
U_G3957: entity G port map(lamdaA => P(3)(829),lamdaB => P(3)(957),s => s(3)(445),lamdaOut => P(2)(957));
U_G3958: entity G port map(lamdaA => P(3)(830),lamdaB => P(3)(958),s => s(3)(446),lamdaOut => P(2)(958));
U_G3959: entity G port map(lamdaA => P(3)(831),lamdaB => P(3)(959),s => s(3)(447),lamdaOut => P(2)(959));
U_G3960: entity G port map(lamdaA => P(3)(832),lamdaB => P(3)(960),s => s(3)(448),lamdaOut => P(2)(960));
U_G3961: entity G port map(lamdaA => P(3)(833),lamdaB => P(3)(961),s => s(3)(449),lamdaOut => P(2)(961));
U_G3962: entity G port map(lamdaA => P(3)(834),lamdaB => P(3)(962),s => s(3)(450),lamdaOut => P(2)(962));
U_G3963: entity G port map(lamdaA => P(3)(835),lamdaB => P(3)(963),s => s(3)(451),lamdaOut => P(2)(963));
U_G3964: entity G port map(lamdaA => P(3)(836),lamdaB => P(3)(964),s => s(3)(452),lamdaOut => P(2)(964));
U_G3965: entity G port map(lamdaA => P(3)(837),lamdaB => P(3)(965),s => s(3)(453),lamdaOut => P(2)(965));
U_G3966: entity G port map(lamdaA => P(3)(838),lamdaB => P(3)(966),s => s(3)(454),lamdaOut => P(2)(966));
U_G3967: entity G port map(lamdaA => P(3)(839),lamdaB => P(3)(967),s => s(3)(455),lamdaOut => P(2)(967));
U_G3968: entity G port map(lamdaA => P(3)(840),lamdaB => P(3)(968),s => s(3)(456),lamdaOut => P(2)(968));
U_G3969: entity G port map(lamdaA => P(3)(841),lamdaB => P(3)(969),s => s(3)(457),lamdaOut => P(2)(969));
U_G3970: entity G port map(lamdaA => P(3)(842),lamdaB => P(3)(970),s => s(3)(458),lamdaOut => P(2)(970));
U_G3971: entity G port map(lamdaA => P(3)(843),lamdaB => P(3)(971),s => s(3)(459),lamdaOut => P(2)(971));
U_G3972: entity G port map(lamdaA => P(3)(844),lamdaB => P(3)(972),s => s(3)(460),lamdaOut => P(2)(972));
U_G3973: entity G port map(lamdaA => P(3)(845),lamdaB => P(3)(973),s => s(3)(461),lamdaOut => P(2)(973));
U_G3974: entity G port map(lamdaA => P(3)(846),lamdaB => P(3)(974),s => s(3)(462),lamdaOut => P(2)(974));
U_G3975: entity G port map(lamdaA => P(3)(847),lamdaB => P(3)(975),s => s(3)(463),lamdaOut => P(2)(975));
U_G3976: entity G port map(lamdaA => P(3)(848),lamdaB => P(3)(976),s => s(3)(464),lamdaOut => P(2)(976));
U_G3977: entity G port map(lamdaA => P(3)(849),lamdaB => P(3)(977),s => s(3)(465),lamdaOut => P(2)(977));
U_G3978: entity G port map(lamdaA => P(3)(850),lamdaB => P(3)(978),s => s(3)(466),lamdaOut => P(2)(978));
U_G3979: entity G port map(lamdaA => P(3)(851),lamdaB => P(3)(979),s => s(3)(467),lamdaOut => P(2)(979));
U_G3980: entity G port map(lamdaA => P(3)(852),lamdaB => P(3)(980),s => s(3)(468),lamdaOut => P(2)(980));
U_G3981: entity G port map(lamdaA => P(3)(853),lamdaB => P(3)(981),s => s(3)(469),lamdaOut => P(2)(981));
U_G3982: entity G port map(lamdaA => P(3)(854),lamdaB => P(3)(982),s => s(3)(470),lamdaOut => P(2)(982));
U_G3983: entity G port map(lamdaA => P(3)(855),lamdaB => P(3)(983),s => s(3)(471),lamdaOut => P(2)(983));
U_G3984: entity G port map(lamdaA => P(3)(856),lamdaB => P(3)(984),s => s(3)(472),lamdaOut => P(2)(984));
U_G3985: entity G port map(lamdaA => P(3)(857),lamdaB => P(3)(985),s => s(3)(473),lamdaOut => P(2)(985));
U_G3986: entity G port map(lamdaA => P(3)(858),lamdaB => P(3)(986),s => s(3)(474),lamdaOut => P(2)(986));
U_G3987: entity G port map(lamdaA => P(3)(859),lamdaB => P(3)(987),s => s(3)(475),lamdaOut => P(2)(987));
U_G3988: entity G port map(lamdaA => P(3)(860),lamdaB => P(3)(988),s => s(3)(476),lamdaOut => P(2)(988));
U_G3989: entity G port map(lamdaA => P(3)(861),lamdaB => P(3)(989),s => s(3)(477),lamdaOut => P(2)(989));
U_G3990: entity G port map(lamdaA => P(3)(862),lamdaB => P(3)(990),s => s(3)(478),lamdaOut => P(2)(990));
U_G3991: entity G port map(lamdaA => P(3)(863),lamdaB => P(3)(991),s => s(3)(479),lamdaOut => P(2)(991));
U_G3992: entity G port map(lamdaA => P(3)(864),lamdaB => P(3)(992),s => s(3)(480),lamdaOut => P(2)(992));
U_G3993: entity G port map(lamdaA => P(3)(865),lamdaB => P(3)(993),s => s(3)(481),lamdaOut => P(2)(993));
U_G3994: entity G port map(lamdaA => P(3)(866),lamdaB => P(3)(994),s => s(3)(482),lamdaOut => P(2)(994));
U_G3995: entity G port map(lamdaA => P(3)(867),lamdaB => P(3)(995),s => s(3)(483),lamdaOut => P(2)(995));
U_G3996: entity G port map(lamdaA => P(3)(868),lamdaB => P(3)(996),s => s(3)(484),lamdaOut => P(2)(996));
U_G3997: entity G port map(lamdaA => P(3)(869),lamdaB => P(3)(997),s => s(3)(485),lamdaOut => P(2)(997));
U_G3998: entity G port map(lamdaA => P(3)(870),lamdaB => P(3)(998),s => s(3)(486),lamdaOut => P(2)(998));
U_G3999: entity G port map(lamdaA => P(3)(871),lamdaB => P(3)(999),s => s(3)(487),lamdaOut => P(2)(999));
U_G31000: entity G port map(lamdaA => P(3)(872),lamdaB => P(3)(1000),s => s(3)(488),lamdaOut => P(2)(1000));
U_G31001: entity G port map(lamdaA => P(3)(873),lamdaB => P(3)(1001),s => s(3)(489),lamdaOut => P(2)(1001));
U_G31002: entity G port map(lamdaA => P(3)(874),lamdaB => P(3)(1002),s => s(3)(490),lamdaOut => P(2)(1002));
U_G31003: entity G port map(lamdaA => P(3)(875),lamdaB => P(3)(1003),s => s(3)(491),lamdaOut => P(2)(1003));
U_G31004: entity G port map(lamdaA => P(3)(876),lamdaB => P(3)(1004),s => s(3)(492),lamdaOut => P(2)(1004));
U_G31005: entity G port map(lamdaA => P(3)(877),lamdaB => P(3)(1005),s => s(3)(493),lamdaOut => P(2)(1005));
U_G31006: entity G port map(lamdaA => P(3)(878),lamdaB => P(3)(1006),s => s(3)(494),lamdaOut => P(2)(1006));
U_G31007: entity G port map(lamdaA => P(3)(879),lamdaB => P(3)(1007),s => s(3)(495),lamdaOut => P(2)(1007));
U_G31008: entity G port map(lamdaA => P(3)(880),lamdaB => P(3)(1008),s => s(3)(496),lamdaOut => P(2)(1008));
U_G31009: entity G port map(lamdaA => P(3)(881),lamdaB => P(3)(1009),s => s(3)(497),lamdaOut => P(2)(1009));
U_G31010: entity G port map(lamdaA => P(3)(882),lamdaB => P(3)(1010),s => s(3)(498),lamdaOut => P(2)(1010));
U_G31011: entity G port map(lamdaA => P(3)(883),lamdaB => P(3)(1011),s => s(3)(499),lamdaOut => P(2)(1011));
U_G31012: entity G port map(lamdaA => P(3)(884),lamdaB => P(3)(1012),s => s(3)(500),lamdaOut => P(2)(1012));
U_G31013: entity G port map(lamdaA => P(3)(885),lamdaB => P(3)(1013),s => s(3)(501),lamdaOut => P(2)(1013));
U_G31014: entity G port map(lamdaA => P(3)(886),lamdaB => P(3)(1014),s => s(3)(502),lamdaOut => P(2)(1014));
U_G31015: entity G port map(lamdaA => P(3)(887),lamdaB => P(3)(1015),s => s(3)(503),lamdaOut => P(2)(1015));
U_G31016: entity G port map(lamdaA => P(3)(888),lamdaB => P(3)(1016),s => s(3)(504),lamdaOut => P(2)(1016));
U_G31017: entity G port map(lamdaA => P(3)(889),lamdaB => P(3)(1017),s => s(3)(505),lamdaOut => P(2)(1017));
U_G31018: entity G port map(lamdaA => P(3)(890),lamdaB => P(3)(1018),s => s(3)(506),lamdaOut => P(2)(1018));
U_G31019: entity G port map(lamdaA => P(3)(891),lamdaB => P(3)(1019),s => s(3)(507),lamdaOut => P(2)(1019));
U_G31020: entity G port map(lamdaA => P(3)(892),lamdaB => P(3)(1020),s => s(3)(508),lamdaOut => P(2)(1020));
U_G31021: entity G port map(lamdaA => P(3)(893),lamdaB => P(3)(1021),s => s(3)(509),lamdaOut => P(2)(1021));
U_G31022: entity G port map(lamdaA => P(3)(894),lamdaB => P(3)(1022),s => s(3)(510),lamdaOut => P(2)(1022));
U_G31023: entity G port map(lamdaA => P(3)(895),lamdaB => P(3)(1023),s => s(3)(511),lamdaOut => P(2)(1023));
-- STAGE 1
U_F20: entity F port map(lamdaA => P(2)(0),lamdaB => P(2)(256),lamdaOut => P(1)(0));
U_F21: entity F port map(lamdaA => P(2)(1),lamdaB => P(2)(257),lamdaOut => P(1)(1));
U_F22: entity F port map(lamdaA => P(2)(2),lamdaB => P(2)(258),lamdaOut => P(1)(2));
U_F23: entity F port map(lamdaA => P(2)(3),lamdaB => P(2)(259),lamdaOut => P(1)(3));
U_F24: entity F port map(lamdaA => P(2)(4),lamdaB => P(2)(260),lamdaOut => P(1)(4));
U_F25: entity F port map(lamdaA => P(2)(5),lamdaB => P(2)(261),lamdaOut => P(1)(5));
U_F26: entity F port map(lamdaA => P(2)(6),lamdaB => P(2)(262),lamdaOut => P(1)(6));
U_F27: entity F port map(lamdaA => P(2)(7),lamdaB => P(2)(263),lamdaOut => P(1)(7));
U_F28: entity F port map(lamdaA => P(2)(8),lamdaB => P(2)(264),lamdaOut => P(1)(8));
U_F29: entity F port map(lamdaA => P(2)(9),lamdaB => P(2)(265),lamdaOut => P(1)(9));
U_F210: entity F port map(lamdaA => P(2)(10),lamdaB => P(2)(266),lamdaOut => P(1)(10));
U_F211: entity F port map(lamdaA => P(2)(11),lamdaB => P(2)(267),lamdaOut => P(1)(11));
U_F212: entity F port map(lamdaA => P(2)(12),lamdaB => P(2)(268),lamdaOut => P(1)(12));
U_F213: entity F port map(lamdaA => P(2)(13),lamdaB => P(2)(269),lamdaOut => P(1)(13));
U_F214: entity F port map(lamdaA => P(2)(14),lamdaB => P(2)(270),lamdaOut => P(1)(14));
U_F215: entity F port map(lamdaA => P(2)(15),lamdaB => P(2)(271),lamdaOut => P(1)(15));
U_F216: entity F port map(lamdaA => P(2)(16),lamdaB => P(2)(272),lamdaOut => P(1)(16));
U_F217: entity F port map(lamdaA => P(2)(17),lamdaB => P(2)(273),lamdaOut => P(1)(17));
U_F218: entity F port map(lamdaA => P(2)(18),lamdaB => P(2)(274),lamdaOut => P(1)(18));
U_F219: entity F port map(lamdaA => P(2)(19),lamdaB => P(2)(275),lamdaOut => P(1)(19));
U_F220: entity F port map(lamdaA => P(2)(20),lamdaB => P(2)(276),lamdaOut => P(1)(20));
U_F221: entity F port map(lamdaA => P(2)(21),lamdaB => P(2)(277),lamdaOut => P(1)(21));
U_F222: entity F port map(lamdaA => P(2)(22),lamdaB => P(2)(278),lamdaOut => P(1)(22));
U_F223: entity F port map(lamdaA => P(2)(23),lamdaB => P(2)(279),lamdaOut => P(1)(23));
U_F224: entity F port map(lamdaA => P(2)(24),lamdaB => P(2)(280),lamdaOut => P(1)(24));
U_F225: entity F port map(lamdaA => P(2)(25),lamdaB => P(2)(281),lamdaOut => P(1)(25));
U_F226: entity F port map(lamdaA => P(2)(26),lamdaB => P(2)(282),lamdaOut => P(1)(26));
U_F227: entity F port map(lamdaA => P(2)(27),lamdaB => P(2)(283),lamdaOut => P(1)(27));
U_F228: entity F port map(lamdaA => P(2)(28),lamdaB => P(2)(284),lamdaOut => P(1)(28));
U_F229: entity F port map(lamdaA => P(2)(29),lamdaB => P(2)(285),lamdaOut => P(1)(29));
U_F230: entity F port map(lamdaA => P(2)(30),lamdaB => P(2)(286),lamdaOut => P(1)(30));
U_F231: entity F port map(lamdaA => P(2)(31),lamdaB => P(2)(287),lamdaOut => P(1)(31));
U_F232: entity F port map(lamdaA => P(2)(32),lamdaB => P(2)(288),lamdaOut => P(1)(32));
U_F233: entity F port map(lamdaA => P(2)(33),lamdaB => P(2)(289),lamdaOut => P(1)(33));
U_F234: entity F port map(lamdaA => P(2)(34),lamdaB => P(2)(290),lamdaOut => P(1)(34));
U_F235: entity F port map(lamdaA => P(2)(35),lamdaB => P(2)(291),lamdaOut => P(1)(35));
U_F236: entity F port map(lamdaA => P(2)(36),lamdaB => P(2)(292),lamdaOut => P(1)(36));
U_F237: entity F port map(lamdaA => P(2)(37),lamdaB => P(2)(293),lamdaOut => P(1)(37));
U_F238: entity F port map(lamdaA => P(2)(38),lamdaB => P(2)(294),lamdaOut => P(1)(38));
U_F239: entity F port map(lamdaA => P(2)(39),lamdaB => P(2)(295),lamdaOut => P(1)(39));
U_F240: entity F port map(lamdaA => P(2)(40),lamdaB => P(2)(296),lamdaOut => P(1)(40));
U_F241: entity F port map(lamdaA => P(2)(41),lamdaB => P(2)(297),lamdaOut => P(1)(41));
U_F242: entity F port map(lamdaA => P(2)(42),lamdaB => P(2)(298),lamdaOut => P(1)(42));
U_F243: entity F port map(lamdaA => P(2)(43),lamdaB => P(2)(299),lamdaOut => P(1)(43));
U_F244: entity F port map(lamdaA => P(2)(44),lamdaB => P(2)(300),lamdaOut => P(1)(44));
U_F245: entity F port map(lamdaA => P(2)(45),lamdaB => P(2)(301),lamdaOut => P(1)(45));
U_F246: entity F port map(lamdaA => P(2)(46),lamdaB => P(2)(302),lamdaOut => P(1)(46));
U_F247: entity F port map(lamdaA => P(2)(47),lamdaB => P(2)(303),lamdaOut => P(1)(47));
U_F248: entity F port map(lamdaA => P(2)(48),lamdaB => P(2)(304),lamdaOut => P(1)(48));
U_F249: entity F port map(lamdaA => P(2)(49),lamdaB => P(2)(305),lamdaOut => P(1)(49));
U_F250: entity F port map(lamdaA => P(2)(50),lamdaB => P(2)(306),lamdaOut => P(1)(50));
U_F251: entity F port map(lamdaA => P(2)(51),lamdaB => P(2)(307),lamdaOut => P(1)(51));
U_F252: entity F port map(lamdaA => P(2)(52),lamdaB => P(2)(308),lamdaOut => P(1)(52));
U_F253: entity F port map(lamdaA => P(2)(53),lamdaB => P(2)(309),lamdaOut => P(1)(53));
U_F254: entity F port map(lamdaA => P(2)(54),lamdaB => P(2)(310),lamdaOut => P(1)(54));
U_F255: entity F port map(lamdaA => P(2)(55),lamdaB => P(2)(311),lamdaOut => P(1)(55));
U_F256: entity F port map(lamdaA => P(2)(56),lamdaB => P(2)(312),lamdaOut => P(1)(56));
U_F257: entity F port map(lamdaA => P(2)(57),lamdaB => P(2)(313),lamdaOut => P(1)(57));
U_F258: entity F port map(lamdaA => P(2)(58),lamdaB => P(2)(314),lamdaOut => P(1)(58));
U_F259: entity F port map(lamdaA => P(2)(59),lamdaB => P(2)(315),lamdaOut => P(1)(59));
U_F260: entity F port map(lamdaA => P(2)(60),lamdaB => P(2)(316),lamdaOut => P(1)(60));
U_F261: entity F port map(lamdaA => P(2)(61),lamdaB => P(2)(317),lamdaOut => P(1)(61));
U_F262: entity F port map(lamdaA => P(2)(62),lamdaB => P(2)(318),lamdaOut => P(1)(62));
U_F263: entity F port map(lamdaA => P(2)(63),lamdaB => P(2)(319),lamdaOut => P(1)(63));
U_F264: entity F port map(lamdaA => P(2)(64),lamdaB => P(2)(320),lamdaOut => P(1)(64));
U_F265: entity F port map(lamdaA => P(2)(65),lamdaB => P(2)(321),lamdaOut => P(1)(65));
U_F266: entity F port map(lamdaA => P(2)(66),lamdaB => P(2)(322),lamdaOut => P(1)(66));
U_F267: entity F port map(lamdaA => P(2)(67),lamdaB => P(2)(323),lamdaOut => P(1)(67));
U_F268: entity F port map(lamdaA => P(2)(68),lamdaB => P(2)(324),lamdaOut => P(1)(68));
U_F269: entity F port map(lamdaA => P(2)(69),lamdaB => P(2)(325),lamdaOut => P(1)(69));
U_F270: entity F port map(lamdaA => P(2)(70),lamdaB => P(2)(326),lamdaOut => P(1)(70));
U_F271: entity F port map(lamdaA => P(2)(71),lamdaB => P(2)(327),lamdaOut => P(1)(71));
U_F272: entity F port map(lamdaA => P(2)(72),lamdaB => P(2)(328),lamdaOut => P(1)(72));
U_F273: entity F port map(lamdaA => P(2)(73),lamdaB => P(2)(329),lamdaOut => P(1)(73));
U_F274: entity F port map(lamdaA => P(2)(74),lamdaB => P(2)(330),lamdaOut => P(1)(74));
U_F275: entity F port map(lamdaA => P(2)(75),lamdaB => P(2)(331),lamdaOut => P(1)(75));
U_F276: entity F port map(lamdaA => P(2)(76),lamdaB => P(2)(332),lamdaOut => P(1)(76));
U_F277: entity F port map(lamdaA => P(2)(77),lamdaB => P(2)(333),lamdaOut => P(1)(77));
U_F278: entity F port map(lamdaA => P(2)(78),lamdaB => P(2)(334),lamdaOut => P(1)(78));
U_F279: entity F port map(lamdaA => P(2)(79),lamdaB => P(2)(335),lamdaOut => P(1)(79));
U_F280: entity F port map(lamdaA => P(2)(80),lamdaB => P(2)(336),lamdaOut => P(1)(80));
U_F281: entity F port map(lamdaA => P(2)(81),lamdaB => P(2)(337),lamdaOut => P(1)(81));
U_F282: entity F port map(lamdaA => P(2)(82),lamdaB => P(2)(338),lamdaOut => P(1)(82));
U_F283: entity F port map(lamdaA => P(2)(83),lamdaB => P(2)(339),lamdaOut => P(1)(83));
U_F284: entity F port map(lamdaA => P(2)(84),lamdaB => P(2)(340),lamdaOut => P(1)(84));
U_F285: entity F port map(lamdaA => P(2)(85),lamdaB => P(2)(341),lamdaOut => P(1)(85));
U_F286: entity F port map(lamdaA => P(2)(86),lamdaB => P(2)(342),lamdaOut => P(1)(86));
U_F287: entity F port map(lamdaA => P(2)(87),lamdaB => P(2)(343),lamdaOut => P(1)(87));
U_F288: entity F port map(lamdaA => P(2)(88),lamdaB => P(2)(344),lamdaOut => P(1)(88));
U_F289: entity F port map(lamdaA => P(2)(89),lamdaB => P(2)(345),lamdaOut => P(1)(89));
U_F290: entity F port map(lamdaA => P(2)(90),lamdaB => P(2)(346),lamdaOut => P(1)(90));
U_F291: entity F port map(lamdaA => P(2)(91),lamdaB => P(2)(347),lamdaOut => P(1)(91));
U_F292: entity F port map(lamdaA => P(2)(92),lamdaB => P(2)(348),lamdaOut => P(1)(92));
U_F293: entity F port map(lamdaA => P(2)(93),lamdaB => P(2)(349),lamdaOut => P(1)(93));
U_F294: entity F port map(lamdaA => P(2)(94),lamdaB => P(2)(350),lamdaOut => P(1)(94));
U_F295: entity F port map(lamdaA => P(2)(95),lamdaB => P(2)(351),lamdaOut => P(1)(95));
U_F296: entity F port map(lamdaA => P(2)(96),lamdaB => P(2)(352),lamdaOut => P(1)(96));
U_F297: entity F port map(lamdaA => P(2)(97),lamdaB => P(2)(353),lamdaOut => P(1)(97));
U_F298: entity F port map(lamdaA => P(2)(98),lamdaB => P(2)(354),lamdaOut => P(1)(98));
U_F299: entity F port map(lamdaA => P(2)(99),lamdaB => P(2)(355),lamdaOut => P(1)(99));
U_F2100: entity F port map(lamdaA => P(2)(100),lamdaB => P(2)(356),lamdaOut => P(1)(100));
U_F2101: entity F port map(lamdaA => P(2)(101),lamdaB => P(2)(357),lamdaOut => P(1)(101));
U_F2102: entity F port map(lamdaA => P(2)(102),lamdaB => P(2)(358),lamdaOut => P(1)(102));
U_F2103: entity F port map(lamdaA => P(2)(103),lamdaB => P(2)(359),lamdaOut => P(1)(103));
U_F2104: entity F port map(lamdaA => P(2)(104),lamdaB => P(2)(360),lamdaOut => P(1)(104));
U_F2105: entity F port map(lamdaA => P(2)(105),lamdaB => P(2)(361),lamdaOut => P(1)(105));
U_F2106: entity F port map(lamdaA => P(2)(106),lamdaB => P(2)(362),lamdaOut => P(1)(106));
U_F2107: entity F port map(lamdaA => P(2)(107),lamdaB => P(2)(363),lamdaOut => P(1)(107));
U_F2108: entity F port map(lamdaA => P(2)(108),lamdaB => P(2)(364),lamdaOut => P(1)(108));
U_F2109: entity F port map(lamdaA => P(2)(109),lamdaB => P(2)(365),lamdaOut => P(1)(109));
U_F2110: entity F port map(lamdaA => P(2)(110),lamdaB => P(2)(366),lamdaOut => P(1)(110));
U_F2111: entity F port map(lamdaA => P(2)(111),lamdaB => P(2)(367),lamdaOut => P(1)(111));
U_F2112: entity F port map(lamdaA => P(2)(112),lamdaB => P(2)(368),lamdaOut => P(1)(112));
U_F2113: entity F port map(lamdaA => P(2)(113),lamdaB => P(2)(369),lamdaOut => P(1)(113));
U_F2114: entity F port map(lamdaA => P(2)(114),lamdaB => P(2)(370),lamdaOut => P(1)(114));
U_F2115: entity F port map(lamdaA => P(2)(115),lamdaB => P(2)(371),lamdaOut => P(1)(115));
U_F2116: entity F port map(lamdaA => P(2)(116),lamdaB => P(2)(372),lamdaOut => P(1)(116));
U_F2117: entity F port map(lamdaA => P(2)(117),lamdaB => P(2)(373),lamdaOut => P(1)(117));
U_F2118: entity F port map(lamdaA => P(2)(118),lamdaB => P(2)(374),lamdaOut => P(1)(118));
U_F2119: entity F port map(lamdaA => P(2)(119),lamdaB => P(2)(375),lamdaOut => P(1)(119));
U_F2120: entity F port map(lamdaA => P(2)(120),lamdaB => P(2)(376),lamdaOut => P(1)(120));
U_F2121: entity F port map(lamdaA => P(2)(121),lamdaB => P(2)(377),lamdaOut => P(1)(121));
U_F2122: entity F port map(lamdaA => P(2)(122),lamdaB => P(2)(378),lamdaOut => P(1)(122));
U_F2123: entity F port map(lamdaA => P(2)(123),lamdaB => P(2)(379),lamdaOut => P(1)(123));
U_F2124: entity F port map(lamdaA => P(2)(124),lamdaB => P(2)(380),lamdaOut => P(1)(124));
U_F2125: entity F port map(lamdaA => P(2)(125),lamdaB => P(2)(381),lamdaOut => P(1)(125));
U_F2126: entity F port map(lamdaA => P(2)(126),lamdaB => P(2)(382),lamdaOut => P(1)(126));
U_F2127: entity F port map(lamdaA => P(2)(127),lamdaB => P(2)(383),lamdaOut => P(1)(127));
U_F2128: entity F port map(lamdaA => P(2)(128),lamdaB => P(2)(384),lamdaOut => P(1)(128));
U_F2129: entity F port map(lamdaA => P(2)(129),lamdaB => P(2)(385),lamdaOut => P(1)(129));
U_F2130: entity F port map(lamdaA => P(2)(130),lamdaB => P(2)(386),lamdaOut => P(1)(130));
U_F2131: entity F port map(lamdaA => P(2)(131),lamdaB => P(2)(387),lamdaOut => P(1)(131));
U_F2132: entity F port map(lamdaA => P(2)(132),lamdaB => P(2)(388),lamdaOut => P(1)(132));
U_F2133: entity F port map(lamdaA => P(2)(133),lamdaB => P(2)(389),lamdaOut => P(1)(133));
U_F2134: entity F port map(lamdaA => P(2)(134),lamdaB => P(2)(390),lamdaOut => P(1)(134));
U_F2135: entity F port map(lamdaA => P(2)(135),lamdaB => P(2)(391),lamdaOut => P(1)(135));
U_F2136: entity F port map(lamdaA => P(2)(136),lamdaB => P(2)(392),lamdaOut => P(1)(136));
U_F2137: entity F port map(lamdaA => P(2)(137),lamdaB => P(2)(393),lamdaOut => P(1)(137));
U_F2138: entity F port map(lamdaA => P(2)(138),lamdaB => P(2)(394),lamdaOut => P(1)(138));
U_F2139: entity F port map(lamdaA => P(2)(139),lamdaB => P(2)(395),lamdaOut => P(1)(139));
U_F2140: entity F port map(lamdaA => P(2)(140),lamdaB => P(2)(396),lamdaOut => P(1)(140));
U_F2141: entity F port map(lamdaA => P(2)(141),lamdaB => P(2)(397),lamdaOut => P(1)(141));
U_F2142: entity F port map(lamdaA => P(2)(142),lamdaB => P(2)(398),lamdaOut => P(1)(142));
U_F2143: entity F port map(lamdaA => P(2)(143),lamdaB => P(2)(399),lamdaOut => P(1)(143));
U_F2144: entity F port map(lamdaA => P(2)(144),lamdaB => P(2)(400),lamdaOut => P(1)(144));
U_F2145: entity F port map(lamdaA => P(2)(145),lamdaB => P(2)(401),lamdaOut => P(1)(145));
U_F2146: entity F port map(lamdaA => P(2)(146),lamdaB => P(2)(402),lamdaOut => P(1)(146));
U_F2147: entity F port map(lamdaA => P(2)(147),lamdaB => P(2)(403),lamdaOut => P(1)(147));
U_F2148: entity F port map(lamdaA => P(2)(148),lamdaB => P(2)(404),lamdaOut => P(1)(148));
U_F2149: entity F port map(lamdaA => P(2)(149),lamdaB => P(2)(405),lamdaOut => P(1)(149));
U_F2150: entity F port map(lamdaA => P(2)(150),lamdaB => P(2)(406),lamdaOut => P(1)(150));
U_F2151: entity F port map(lamdaA => P(2)(151),lamdaB => P(2)(407),lamdaOut => P(1)(151));
U_F2152: entity F port map(lamdaA => P(2)(152),lamdaB => P(2)(408),lamdaOut => P(1)(152));
U_F2153: entity F port map(lamdaA => P(2)(153),lamdaB => P(2)(409),lamdaOut => P(1)(153));
U_F2154: entity F port map(lamdaA => P(2)(154),lamdaB => P(2)(410),lamdaOut => P(1)(154));
U_F2155: entity F port map(lamdaA => P(2)(155),lamdaB => P(2)(411),lamdaOut => P(1)(155));
U_F2156: entity F port map(lamdaA => P(2)(156),lamdaB => P(2)(412),lamdaOut => P(1)(156));
U_F2157: entity F port map(lamdaA => P(2)(157),lamdaB => P(2)(413),lamdaOut => P(1)(157));
U_F2158: entity F port map(lamdaA => P(2)(158),lamdaB => P(2)(414),lamdaOut => P(1)(158));
U_F2159: entity F port map(lamdaA => P(2)(159),lamdaB => P(2)(415),lamdaOut => P(1)(159));
U_F2160: entity F port map(lamdaA => P(2)(160),lamdaB => P(2)(416),lamdaOut => P(1)(160));
U_F2161: entity F port map(lamdaA => P(2)(161),lamdaB => P(2)(417),lamdaOut => P(1)(161));
U_F2162: entity F port map(lamdaA => P(2)(162),lamdaB => P(2)(418),lamdaOut => P(1)(162));
U_F2163: entity F port map(lamdaA => P(2)(163),lamdaB => P(2)(419),lamdaOut => P(1)(163));
U_F2164: entity F port map(lamdaA => P(2)(164),lamdaB => P(2)(420),lamdaOut => P(1)(164));
U_F2165: entity F port map(lamdaA => P(2)(165),lamdaB => P(2)(421),lamdaOut => P(1)(165));
U_F2166: entity F port map(lamdaA => P(2)(166),lamdaB => P(2)(422),lamdaOut => P(1)(166));
U_F2167: entity F port map(lamdaA => P(2)(167),lamdaB => P(2)(423),lamdaOut => P(1)(167));
U_F2168: entity F port map(lamdaA => P(2)(168),lamdaB => P(2)(424),lamdaOut => P(1)(168));
U_F2169: entity F port map(lamdaA => P(2)(169),lamdaB => P(2)(425),lamdaOut => P(1)(169));
U_F2170: entity F port map(lamdaA => P(2)(170),lamdaB => P(2)(426),lamdaOut => P(1)(170));
U_F2171: entity F port map(lamdaA => P(2)(171),lamdaB => P(2)(427),lamdaOut => P(1)(171));
U_F2172: entity F port map(lamdaA => P(2)(172),lamdaB => P(2)(428),lamdaOut => P(1)(172));
U_F2173: entity F port map(lamdaA => P(2)(173),lamdaB => P(2)(429),lamdaOut => P(1)(173));
U_F2174: entity F port map(lamdaA => P(2)(174),lamdaB => P(2)(430),lamdaOut => P(1)(174));
U_F2175: entity F port map(lamdaA => P(2)(175),lamdaB => P(2)(431),lamdaOut => P(1)(175));
U_F2176: entity F port map(lamdaA => P(2)(176),lamdaB => P(2)(432),lamdaOut => P(1)(176));
U_F2177: entity F port map(lamdaA => P(2)(177),lamdaB => P(2)(433),lamdaOut => P(1)(177));
U_F2178: entity F port map(lamdaA => P(2)(178),lamdaB => P(2)(434),lamdaOut => P(1)(178));
U_F2179: entity F port map(lamdaA => P(2)(179),lamdaB => P(2)(435),lamdaOut => P(1)(179));
U_F2180: entity F port map(lamdaA => P(2)(180),lamdaB => P(2)(436),lamdaOut => P(1)(180));
U_F2181: entity F port map(lamdaA => P(2)(181),lamdaB => P(2)(437),lamdaOut => P(1)(181));
U_F2182: entity F port map(lamdaA => P(2)(182),lamdaB => P(2)(438),lamdaOut => P(1)(182));
U_F2183: entity F port map(lamdaA => P(2)(183),lamdaB => P(2)(439),lamdaOut => P(1)(183));
U_F2184: entity F port map(lamdaA => P(2)(184),lamdaB => P(2)(440),lamdaOut => P(1)(184));
U_F2185: entity F port map(lamdaA => P(2)(185),lamdaB => P(2)(441),lamdaOut => P(1)(185));
U_F2186: entity F port map(lamdaA => P(2)(186),lamdaB => P(2)(442),lamdaOut => P(1)(186));
U_F2187: entity F port map(lamdaA => P(2)(187),lamdaB => P(2)(443),lamdaOut => P(1)(187));
U_F2188: entity F port map(lamdaA => P(2)(188),lamdaB => P(2)(444),lamdaOut => P(1)(188));
U_F2189: entity F port map(lamdaA => P(2)(189),lamdaB => P(2)(445),lamdaOut => P(1)(189));
U_F2190: entity F port map(lamdaA => P(2)(190),lamdaB => P(2)(446),lamdaOut => P(1)(190));
U_F2191: entity F port map(lamdaA => P(2)(191),lamdaB => P(2)(447),lamdaOut => P(1)(191));
U_F2192: entity F port map(lamdaA => P(2)(192),lamdaB => P(2)(448),lamdaOut => P(1)(192));
U_F2193: entity F port map(lamdaA => P(2)(193),lamdaB => P(2)(449),lamdaOut => P(1)(193));
U_F2194: entity F port map(lamdaA => P(2)(194),lamdaB => P(2)(450),lamdaOut => P(1)(194));
U_F2195: entity F port map(lamdaA => P(2)(195),lamdaB => P(2)(451),lamdaOut => P(1)(195));
U_F2196: entity F port map(lamdaA => P(2)(196),lamdaB => P(2)(452),lamdaOut => P(1)(196));
U_F2197: entity F port map(lamdaA => P(2)(197),lamdaB => P(2)(453),lamdaOut => P(1)(197));
U_F2198: entity F port map(lamdaA => P(2)(198),lamdaB => P(2)(454),lamdaOut => P(1)(198));
U_F2199: entity F port map(lamdaA => P(2)(199),lamdaB => P(2)(455),lamdaOut => P(1)(199));
U_F2200: entity F port map(lamdaA => P(2)(200),lamdaB => P(2)(456),lamdaOut => P(1)(200));
U_F2201: entity F port map(lamdaA => P(2)(201),lamdaB => P(2)(457),lamdaOut => P(1)(201));
U_F2202: entity F port map(lamdaA => P(2)(202),lamdaB => P(2)(458),lamdaOut => P(1)(202));
U_F2203: entity F port map(lamdaA => P(2)(203),lamdaB => P(2)(459),lamdaOut => P(1)(203));
U_F2204: entity F port map(lamdaA => P(2)(204),lamdaB => P(2)(460),lamdaOut => P(1)(204));
U_F2205: entity F port map(lamdaA => P(2)(205),lamdaB => P(2)(461),lamdaOut => P(1)(205));
U_F2206: entity F port map(lamdaA => P(2)(206),lamdaB => P(2)(462),lamdaOut => P(1)(206));
U_F2207: entity F port map(lamdaA => P(2)(207),lamdaB => P(2)(463),lamdaOut => P(1)(207));
U_F2208: entity F port map(lamdaA => P(2)(208),lamdaB => P(2)(464),lamdaOut => P(1)(208));
U_F2209: entity F port map(lamdaA => P(2)(209),lamdaB => P(2)(465),lamdaOut => P(1)(209));
U_F2210: entity F port map(lamdaA => P(2)(210),lamdaB => P(2)(466),lamdaOut => P(1)(210));
U_F2211: entity F port map(lamdaA => P(2)(211),lamdaB => P(2)(467),lamdaOut => P(1)(211));
U_F2212: entity F port map(lamdaA => P(2)(212),lamdaB => P(2)(468),lamdaOut => P(1)(212));
U_F2213: entity F port map(lamdaA => P(2)(213),lamdaB => P(2)(469),lamdaOut => P(1)(213));
U_F2214: entity F port map(lamdaA => P(2)(214),lamdaB => P(2)(470),lamdaOut => P(1)(214));
U_F2215: entity F port map(lamdaA => P(2)(215),lamdaB => P(2)(471),lamdaOut => P(1)(215));
U_F2216: entity F port map(lamdaA => P(2)(216),lamdaB => P(2)(472),lamdaOut => P(1)(216));
U_F2217: entity F port map(lamdaA => P(2)(217),lamdaB => P(2)(473),lamdaOut => P(1)(217));
U_F2218: entity F port map(lamdaA => P(2)(218),lamdaB => P(2)(474),lamdaOut => P(1)(218));
U_F2219: entity F port map(lamdaA => P(2)(219),lamdaB => P(2)(475),lamdaOut => P(1)(219));
U_F2220: entity F port map(lamdaA => P(2)(220),lamdaB => P(2)(476),lamdaOut => P(1)(220));
U_F2221: entity F port map(lamdaA => P(2)(221),lamdaB => P(2)(477),lamdaOut => P(1)(221));
U_F2222: entity F port map(lamdaA => P(2)(222),lamdaB => P(2)(478),lamdaOut => P(1)(222));
U_F2223: entity F port map(lamdaA => P(2)(223),lamdaB => P(2)(479),lamdaOut => P(1)(223));
U_F2224: entity F port map(lamdaA => P(2)(224),lamdaB => P(2)(480),lamdaOut => P(1)(224));
U_F2225: entity F port map(lamdaA => P(2)(225),lamdaB => P(2)(481),lamdaOut => P(1)(225));
U_F2226: entity F port map(lamdaA => P(2)(226),lamdaB => P(2)(482),lamdaOut => P(1)(226));
U_F2227: entity F port map(lamdaA => P(2)(227),lamdaB => P(2)(483),lamdaOut => P(1)(227));
U_F2228: entity F port map(lamdaA => P(2)(228),lamdaB => P(2)(484),lamdaOut => P(1)(228));
U_F2229: entity F port map(lamdaA => P(2)(229),lamdaB => P(2)(485),lamdaOut => P(1)(229));
U_F2230: entity F port map(lamdaA => P(2)(230),lamdaB => P(2)(486),lamdaOut => P(1)(230));
U_F2231: entity F port map(lamdaA => P(2)(231),lamdaB => P(2)(487),lamdaOut => P(1)(231));
U_F2232: entity F port map(lamdaA => P(2)(232),lamdaB => P(2)(488),lamdaOut => P(1)(232));
U_F2233: entity F port map(lamdaA => P(2)(233),lamdaB => P(2)(489),lamdaOut => P(1)(233));
U_F2234: entity F port map(lamdaA => P(2)(234),lamdaB => P(2)(490),lamdaOut => P(1)(234));
U_F2235: entity F port map(lamdaA => P(2)(235),lamdaB => P(2)(491),lamdaOut => P(1)(235));
U_F2236: entity F port map(lamdaA => P(2)(236),lamdaB => P(2)(492),lamdaOut => P(1)(236));
U_F2237: entity F port map(lamdaA => P(2)(237),lamdaB => P(2)(493),lamdaOut => P(1)(237));
U_F2238: entity F port map(lamdaA => P(2)(238),lamdaB => P(2)(494),lamdaOut => P(1)(238));
U_F2239: entity F port map(lamdaA => P(2)(239),lamdaB => P(2)(495),lamdaOut => P(1)(239));
U_F2240: entity F port map(lamdaA => P(2)(240),lamdaB => P(2)(496),lamdaOut => P(1)(240));
U_F2241: entity F port map(lamdaA => P(2)(241),lamdaB => P(2)(497),lamdaOut => P(1)(241));
U_F2242: entity F port map(lamdaA => P(2)(242),lamdaB => P(2)(498),lamdaOut => P(1)(242));
U_F2243: entity F port map(lamdaA => P(2)(243),lamdaB => P(2)(499),lamdaOut => P(1)(243));
U_F2244: entity F port map(lamdaA => P(2)(244),lamdaB => P(2)(500),lamdaOut => P(1)(244));
U_F2245: entity F port map(lamdaA => P(2)(245),lamdaB => P(2)(501),lamdaOut => P(1)(245));
U_F2246: entity F port map(lamdaA => P(2)(246),lamdaB => P(2)(502),lamdaOut => P(1)(246));
U_F2247: entity F port map(lamdaA => P(2)(247),lamdaB => P(2)(503),lamdaOut => P(1)(247));
U_F2248: entity F port map(lamdaA => P(2)(248),lamdaB => P(2)(504),lamdaOut => P(1)(248));
U_F2249: entity F port map(lamdaA => P(2)(249),lamdaB => P(2)(505),lamdaOut => P(1)(249));
U_F2250: entity F port map(lamdaA => P(2)(250),lamdaB => P(2)(506),lamdaOut => P(1)(250));
U_F2251: entity F port map(lamdaA => P(2)(251),lamdaB => P(2)(507),lamdaOut => P(1)(251));
U_F2252: entity F port map(lamdaA => P(2)(252),lamdaB => P(2)(508),lamdaOut => P(1)(252));
U_F2253: entity F port map(lamdaA => P(2)(253),lamdaB => P(2)(509),lamdaOut => P(1)(253));
U_F2254: entity F port map(lamdaA => P(2)(254),lamdaB => P(2)(510),lamdaOut => P(1)(254));
U_F2255: entity F port map(lamdaA => P(2)(255),lamdaB => P(2)(511),lamdaOut => P(1)(255));
U_G2256: entity G port map(lamdaA => P(2)(0),lamdaB => P(2)(256),s => s(2)(0),lamdaOut => P(1)(256));
U_G2257: entity G port map(lamdaA => P(2)(1),lamdaB => P(2)(257),s => s(2)(1),lamdaOut => P(1)(257));
U_G2258: entity G port map(lamdaA => P(2)(2),lamdaB => P(2)(258),s => s(2)(2),lamdaOut => P(1)(258));
U_G2259: entity G port map(lamdaA => P(2)(3),lamdaB => P(2)(259),s => s(2)(3),lamdaOut => P(1)(259));
U_G2260: entity G port map(lamdaA => P(2)(4),lamdaB => P(2)(260),s => s(2)(4),lamdaOut => P(1)(260));
U_G2261: entity G port map(lamdaA => P(2)(5),lamdaB => P(2)(261),s => s(2)(5),lamdaOut => P(1)(261));
U_G2262: entity G port map(lamdaA => P(2)(6),lamdaB => P(2)(262),s => s(2)(6),lamdaOut => P(1)(262));
U_G2263: entity G port map(lamdaA => P(2)(7),lamdaB => P(2)(263),s => s(2)(7),lamdaOut => P(1)(263));
U_G2264: entity G port map(lamdaA => P(2)(8),lamdaB => P(2)(264),s => s(2)(8),lamdaOut => P(1)(264));
U_G2265: entity G port map(lamdaA => P(2)(9),lamdaB => P(2)(265),s => s(2)(9),lamdaOut => P(1)(265));
U_G2266: entity G port map(lamdaA => P(2)(10),lamdaB => P(2)(266),s => s(2)(10),lamdaOut => P(1)(266));
U_G2267: entity G port map(lamdaA => P(2)(11),lamdaB => P(2)(267),s => s(2)(11),lamdaOut => P(1)(267));
U_G2268: entity G port map(lamdaA => P(2)(12),lamdaB => P(2)(268),s => s(2)(12),lamdaOut => P(1)(268));
U_G2269: entity G port map(lamdaA => P(2)(13),lamdaB => P(2)(269),s => s(2)(13),lamdaOut => P(1)(269));
U_G2270: entity G port map(lamdaA => P(2)(14),lamdaB => P(2)(270),s => s(2)(14),lamdaOut => P(1)(270));
U_G2271: entity G port map(lamdaA => P(2)(15),lamdaB => P(2)(271),s => s(2)(15),lamdaOut => P(1)(271));
U_G2272: entity G port map(lamdaA => P(2)(16),lamdaB => P(2)(272),s => s(2)(16),lamdaOut => P(1)(272));
U_G2273: entity G port map(lamdaA => P(2)(17),lamdaB => P(2)(273),s => s(2)(17),lamdaOut => P(1)(273));
U_G2274: entity G port map(lamdaA => P(2)(18),lamdaB => P(2)(274),s => s(2)(18),lamdaOut => P(1)(274));
U_G2275: entity G port map(lamdaA => P(2)(19),lamdaB => P(2)(275),s => s(2)(19),lamdaOut => P(1)(275));
U_G2276: entity G port map(lamdaA => P(2)(20),lamdaB => P(2)(276),s => s(2)(20),lamdaOut => P(1)(276));
U_G2277: entity G port map(lamdaA => P(2)(21),lamdaB => P(2)(277),s => s(2)(21),lamdaOut => P(1)(277));
U_G2278: entity G port map(lamdaA => P(2)(22),lamdaB => P(2)(278),s => s(2)(22),lamdaOut => P(1)(278));
U_G2279: entity G port map(lamdaA => P(2)(23),lamdaB => P(2)(279),s => s(2)(23),lamdaOut => P(1)(279));
U_G2280: entity G port map(lamdaA => P(2)(24),lamdaB => P(2)(280),s => s(2)(24),lamdaOut => P(1)(280));
U_G2281: entity G port map(lamdaA => P(2)(25),lamdaB => P(2)(281),s => s(2)(25),lamdaOut => P(1)(281));
U_G2282: entity G port map(lamdaA => P(2)(26),lamdaB => P(2)(282),s => s(2)(26),lamdaOut => P(1)(282));
U_G2283: entity G port map(lamdaA => P(2)(27),lamdaB => P(2)(283),s => s(2)(27),lamdaOut => P(1)(283));
U_G2284: entity G port map(lamdaA => P(2)(28),lamdaB => P(2)(284),s => s(2)(28),lamdaOut => P(1)(284));
U_G2285: entity G port map(lamdaA => P(2)(29),lamdaB => P(2)(285),s => s(2)(29),lamdaOut => P(1)(285));
U_G2286: entity G port map(lamdaA => P(2)(30),lamdaB => P(2)(286),s => s(2)(30),lamdaOut => P(1)(286));
U_G2287: entity G port map(lamdaA => P(2)(31),lamdaB => P(2)(287),s => s(2)(31),lamdaOut => P(1)(287));
U_G2288: entity G port map(lamdaA => P(2)(32),lamdaB => P(2)(288),s => s(2)(32),lamdaOut => P(1)(288));
U_G2289: entity G port map(lamdaA => P(2)(33),lamdaB => P(2)(289),s => s(2)(33),lamdaOut => P(1)(289));
U_G2290: entity G port map(lamdaA => P(2)(34),lamdaB => P(2)(290),s => s(2)(34),lamdaOut => P(1)(290));
U_G2291: entity G port map(lamdaA => P(2)(35),lamdaB => P(2)(291),s => s(2)(35),lamdaOut => P(1)(291));
U_G2292: entity G port map(lamdaA => P(2)(36),lamdaB => P(2)(292),s => s(2)(36),lamdaOut => P(1)(292));
U_G2293: entity G port map(lamdaA => P(2)(37),lamdaB => P(2)(293),s => s(2)(37),lamdaOut => P(1)(293));
U_G2294: entity G port map(lamdaA => P(2)(38),lamdaB => P(2)(294),s => s(2)(38),lamdaOut => P(1)(294));
U_G2295: entity G port map(lamdaA => P(2)(39),lamdaB => P(2)(295),s => s(2)(39),lamdaOut => P(1)(295));
U_G2296: entity G port map(lamdaA => P(2)(40),lamdaB => P(2)(296),s => s(2)(40),lamdaOut => P(1)(296));
U_G2297: entity G port map(lamdaA => P(2)(41),lamdaB => P(2)(297),s => s(2)(41),lamdaOut => P(1)(297));
U_G2298: entity G port map(lamdaA => P(2)(42),lamdaB => P(2)(298),s => s(2)(42),lamdaOut => P(1)(298));
U_G2299: entity G port map(lamdaA => P(2)(43),lamdaB => P(2)(299),s => s(2)(43),lamdaOut => P(1)(299));
U_G2300: entity G port map(lamdaA => P(2)(44),lamdaB => P(2)(300),s => s(2)(44),lamdaOut => P(1)(300));
U_G2301: entity G port map(lamdaA => P(2)(45),lamdaB => P(2)(301),s => s(2)(45),lamdaOut => P(1)(301));
U_G2302: entity G port map(lamdaA => P(2)(46),lamdaB => P(2)(302),s => s(2)(46),lamdaOut => P(1)(302));
U_G2303: entity G port map(lamdaA => P(2)(47),lamdaB => P(2)(303),s => s(2)(47),lamdaOut => P(1)(303));
U_G2304: entity G port map(lamdaA => P(2)(48),lamdaB => P(2)(304),s => s(2)(48),lamdaOut => P(1)(304));
U_G2305: entity G port map(lamdaA => P(2)(49),lamdaB => P(2)(305),s => s(2)(49),lamdaOut => P(1)(305));
U_G2306: entity G port map(lamdaA => P(2)(50),lamdaB => P(2)(306),s => s(2)(50),lamdaOut => P(1)(306));
U_G2307: entity G port map(lamdaA => P(2)(51),lamdaB => P(2)(307),s => s(2)(51),lamdaOut => P(1)(307));
U_G2308: entity G port map(lamdaA => P(2)(52),lamdaB => P(2)(308),s => s(2)(52),lamdaOut => P(1)(308));
U_G2309: entity G port map(lamdaA => P(2)(53),lamdaB => P(2)(309),s => s(2)(53),lamdaOut => P(1)(309));
U_G2310: entity G port map(lamdaA => P(2)(54),lamdaB => P(2)(310),s => s(2)(54),lamdaOut => P(1)(310));
U_G2311: entity G port map(lamdaA => P(2)(55),lamdaB => P(2)(311),s => s(2)(55),lamdaOut => P(1)(311));
U_G2312: entity G port map(lamdaA => P(2)(56),lamdaB => P(2)(312),s => s(2)(56),lamdaOut => P(1)(312));
U_G2313: entity G port map(lamdaA => P(2)(57),lamdaB => P(2)(313),s => s(2)(57),lamdaOut => P(1)(313));
U_G2314: entity G port map(lamdaA => P(2)(58),lamdaB => P(2)(314),s => s(2)(58),lamdaOut => P(1)(314));
U_G2315: entity G port map(lamdaA => P(2)(59),lamdaB => P(2)(315),s => s(2)(59),lamdaOut => P(1)(315));
U_G2316: entity G port map(lamdaA => P(2)(60),lamdaB => P(2)(316),s => s(2)(60),lamdaOut => P(1)(316));
U_G2317: entity G port map(lamdaA => P(2)(61),lamdaB => P(2)(317),s => s(2)(61),lamdaOut => P(1)(317));
U_G2318: entity G port map(lamdaA => P(2)(62),lamdaB => P(2)(318),s => s(2)(62),lamdaOut => P(1)(318));
U_G2319: entity G port map(lamdaA => P(2)(63),lamdaB => P(2)(319),s => s(2)(63),lamdaOut => P(1)(319));
U_G2320: entity G port map(lamdaA => P(2)(64),lamdaB => P(2)(320),s => s(2)(64),lamdaOut => P(1)(320));
U_G2321: entity G port map(lamdaA => P(2)(65),lamdaB => P(2)(321),s => s(2)(65),lamdaOut => P(1)(321));
U_G2322: entity G port map(lamdaA => P(2)(66),lamdaB => P(2)(322),s => s(2)(66),lamdaOut => P(1)(322));
U_G2323: entity G port map(lamdaA => P(2)(67),lamdaB => P(2)(323),s => s(2)(67),lamdaOut => P(1)(323));
U_G2324: entity G port map(lamdaA => P(2)(68),lamdaB => P(2)(324),s => s(2)(68),lamdaOut => P(1)(324));
U_G2325: entity G port map(lamdaA => P(2)(69),lamdaB => P(2)(325),s => s(2)(69),lamdaOut => P(1)(325));
U_G2326: entity G port map(lamdaA => P(2)(70),lamdaB => P(2)(326),s => s(2)(70),lamdaOut => P(1)(326));
U_G2327: entity G port map(lamdaA => P(2)(71),lamdaB => P(2)(327),s => s(2)(71),lamdaOut => P(1)(327));
U_G2328: entity G port map(lamdaA => P(2)(72),lamdaB => P(2)(328),s => s(2)(72),lamdaOut => P(1)(328));
U_G2329: entity G port map(lamdaA => P(2)(73),lamdaB => P(2)(329),s => s(2)(73),lamdaOut => P(1)(329));
U_G2330: entity G port map(lamdaA => P(2)(74),lamdaB => P(2)(330),s => s(2)(74),lamdaOut => P(1)(330));
U_G2331: entity G port map(lamdaA => P(2)(75),lamdaB => P(2)(331),s => s(2)(75),lamdaOut => P(1)(331));
U_G2332: entity G port map(lamdaA => P(2)(76),lamdaB => P(2)(332),s => s(2)(76),lamdaOut => P(1)(332));
U_G2333: entity G port map(lamdaA => P(2)(77),lamdaB => P(2)(333),s => s(2)(77),lamdaOut => P(1)(333));
U_G2334: entity G port map(lamdaA => P(2)(78),lamdaB => P(2)(334),s => s(2)(78),lamdaOut => P(1)(334));
U_G2335: entity G port map(lamdaA => P(2)(79),lamdaB => P(2)(335),s => s(2)(79),lamdaOut => P(1)(335));
U_G2336: entity G port map(lamdaA => P(2)(80),lamdaB => P(2)(336),s => s(2)(80),lamdaOut => P(1)(336));
U_G2337: entity G port map(lamdaA => P(2)(81),lamdaB => P(2)(337),s => s(2)(81),lamdaOut => P(1)(337));
U_G2338: entity G port map(lamdaA => P(2)(82),lamdaB => P(2)(338),s => s(2)(82),lamdaOut => P(1)(338));
U_G2339: entity G port map(lamdaA => P(2)(83),lamdaB => P(2)(339),s => s(2)(83),lamdaOut => P(1)(339));
U_G2340: entity G port map(lamdaA => P(2)(84),lamdaB => P(2)(340),s => s(2)(84),lamdaOut => P(1)(340));
U_G2341: entity G port map(lamdaA => P(2)(85),lamdaB => P(2)(341),s => s(2)(85),lamdaOut => P(1)(341));
U_G2342: entity G port map(lamdaA => P(2)(86),lamdaB => P(2)(342),s => s(2)(86),lamdaOut => P(1)(342));
U_G2343: entity G port map(lamdaA => P(2)(87),lamdaB => P(2)(343),s => s(2)(87),lamdaOut => P(1)(343));
U_G2344: entity G port map(lamdaA => P(2)(88),lamdaB => P(2)(344),s => s(2)(88),lamdaOut => P(1)(344));
U_G2345: entity G port map(lamdaA => P(2)(89),lamdaB => P(2)(345),s => s(2)(89),lamdaOut => P(1)(345));
U_G2346: entity G port map(lamdaA => P(2)(90),lamdaB => P(2)(346),s => s(2)(90),lamdaOut => P(1)(346));
U_G2347: entity G port map(lamdaA => P(2)(91),lamdaB => P(2)(347),s => s(2)(91),lamdaOut => P(1)(347));
U_G2348: entity G port map(lamdaA => P(2)(92),lamdaB => P(2)(348),s => s(2)(92),lamdaOut => P(1)(348));
U_G2349: entity G port map(lamdaA => P(2)(93),lamdaB => P(2)(349),s => s(2)(93),lamdaOut => P(1)(349));
U_G2350: entity G port map(lamdaA => P(2)(94),lamdaB => P(2)(350),s => s(2)(94),lamdaOut => P(1)(350));
U_G2351: entity G port map(lamdaA => P(2)(95),lamdaB => P(2)(351),s => s(2)(95),lamdaOut => P(1)(351));
U_G2352: entity G port map(lamdaA => P(2)(96),lamdaB => P(2)(352),s => s(2)(96),lamdaOut => P(1)(352));
U_G2353: entity G port map(lamdaA => P(2)(97),lamdaB => P(2)(353),s => s(2)(97),lamdaOut => P(1)(353));
U_G2354: entity G port map(lamdaA => P(2)(98),lamdaB => P(2)(354),s => s(2)(98),lamdaOut => P(1)(354));
U_G2355: entity G port map(lamdaA => P(2)(99),lamdaB => P(2)(355),s => s(2)(99),lamdaOut => P(1)(355));
U_G2356: entity G port map(lamdaA => P(2)(100),lamdaB => P(2)(356),s => s(2)(100),lamdaOut => P(1)(356));
U_G2357: entity G port map(lamdaA => P(2)(101),lamdaB => P(2)(357),s => s(2)(101),lamdaOut => P(1)(357));
U_G2358: entity G port map(lamdaA => P(2)(102),lamdaB => P(2)(358),s => s(2)(102),lamdaOut => P(1)(358));
U_G2359: entity G port map(lamdaA => P(2)(103),lamdaB => P(2)(359),s => s(2)(103),lamdaOut => P(1)(359));
U_G2360: entity G port map(lamdaA => P(2)(104),lamdaB => P(2)(360),s => s(2)(104),lamdaOut => P(1)(360));
U_G2361: entity G port map(lamdaA => P(2)(105),lamdaB => P(2)(361),s => s(2)(105),lamdaOut => P(1)(361));
U_G2362: entity G port map(lamdaA => P(2)(106),lamdaB => P(2)(362),s => s(2)(106),lamdaOut => P(1)(362));
U_G2363: entity G port map(lamdaA => P(2)(107),lamdaB => P(2)(363),s => s(2)(107),lamdaOut => P(1)(363));
U_G2364: entity G port map(lamdaA => P(2)(108),lamdaB => P(2)(364),s => s(2)(108),lamdaOut => P(1)(364));
U_G2365: entity G port map(lamdaA => P(2)(109),lamdaB => P(2)(365),s => s(2)(109),lamdaOut => P(1)(365));
U_G2366: entity G port map(lamdaA => P(2)(110),lamdaB => P(2)(366),s => s(2)(110),lamdaOut => P(1)(366));
U_G2367: entity G port map(lamdaA => P(2)(111),lamdaB => P(2)(367),s => s(2)(111),lamdaOut => P(1)(367));
U_G2368: entity G port map(lamdaA => P(2)(112),lamdaB => P(2)(368),s => s(2)(112),lamdaOut => P(1)(368));
U_G2369: entity G port map(lamdaA => P(2)(113),lamdaB => P(2)(369),s => s(2)(113),lamdaOut => P(1)(369));
U_G2370: entity G port map(lamdaA => P(2)(114),lamdaB => P(2)(370),s => s(2)(114),lamdaOut => P(1)(370));
U_G2371: entity G port map(lamdaA => P(2)(115),lamdaB => P(2)(371),s => s(2)(115),lamdaOut => P(1)(371));
U_G2372: entity G port map(lamdaA => P(2)(116),lamdaB => P(2)(372),s => s(2)(116),lamdaOut => P(1)(372));
U_G2373: entity G port map(lamdaA => P(2)(117),lamdaB => P(2)(373),s => s(2)(117),lamdaOut => P(1)(373));
U_G2374: entity G port map(lamdaA => P(2)(118),lamdaB => P(2)(374),s => s(2)(118),lamdaOut => P(1)(374));
U_G2375: entity G port map(lamdaA => P(2)(119),lamdaB => P(2)(375),s => s(2)(119),lamdaOut => P(1)(375));
U_G2376: entity G port map(lamdaA => P(2)(120),lamdaB => P(2)(376),s => s(2)(120),lamdaOut => P(1)(376));
U_G2377: entity G port map(lamdaA => P(2)(121),lamdaB => P(2)(377),s => s(2)(121),lamdaOut => P(1)(377));
U_G2378: entity G port map(lamdaA => P(2)(122),lamdaB => P(2)(378),s => s(2)(122),lamdaOut => P(1)(378));
U_G2379: entity G port map(lamdaA => P(2)(123),lamdaB => P(2)(379),s => s(2)(123),lamdaOut => P(1)(379));
U_G2380: entity G port map(lamdaA => P(2)(124),lamdaB => P(2)(380),s => s(2)(124),lamdaOut => P(1)(380));
U_G2381: entity G port map(lamdaA => P(2)(125),lamdaB => P(2)(381),s => s(2)(125),lamdaOut => P(1)(381));
U_G2382: entity G port map(lamdaA => P(2)(126),lamdaB => P(2)(382),s => s(2)(126),lamdaOut => P(1)(382));
U_G2383: entity G port map(lamdaA => P(2)(127),lamdaB => P(2)(383),s => s(2)(127),lamdaOut => P(1)(383));
U_G2384: entity G port map(lamdaA => P(2)(128),lamdaB => P(2)(384),s => s(2)(128),lamdaOut => P(1)(384));
U_G2385: entity G port map(lamdaA => P(2)(129),lamdaB => P(2)(385),s => s(2)(129),lamdaOut => P(1)(385));
U_G2386: entity G port map(lamdaA => P(2)(130),lamdaB => P(2)(386),s => s(2)(130),lamdaOut => P(1)(386));
U_G2387: entity G port map(lamdaA => P(2)(131),lamdaB => P(2)(387),s => s(2)(131),lamdaOut => P(1)(387));
U_G2388: entity G port map(lamdaA => P(2)(132),lamdaB => P(2)(388),s => s(2)(132),lamdaOut => P(1)(388));
U_G2389: entity G port map(lamdaA => P(2)(133),lamdaB => P(2)(389),s => s(2)(133),lamdaOut => P(1)(389));
U_G2390: entity G port map(lamdaA => P(2)(134),lamdaB => P(2)(390),s => s(2)(134),lamdaOut => P(1)(390));
U_G2391: entity G port map(lamdaA => P(2)(135),lamdaB => P(2)(391),s => s(2)(135),lamdaOut => P(1)(391));
U_G2392: entity G port map(lamdaA => P(2)(136),lamdaB => P(2)(392),s => s(2)(136),lamdaOut => P(1)(392));
U_G2393: entity G port map(lamdaA => P(2)(137),lamdaB => P(2)(393),s => s(2)(137),lamdaOut => P(1)(393));
U_G2394: entity G port map(lamdaA => P(2)(138),lamdaB => P(2)(394),s => s(2)(138),lamdaOut => P(1)(394));
U_G2395: entity G port map(lamdaA => P(2)(139),lamdaB => P(2)(395),s => s(2)(139),lamdaOut => P(1)(395));
U_G2396: entity G port map(lamdaA => P(2)(140),lamdaB => P(2)(396),s => s(2)(140),lamdaOut => P(1)(396));
U_G2397: entity G port map(lamdaA => P(2)(141),lamdaB => P(2)(397),s => s(2)(141),lamdaOut => P(1)(397));
U_G2398: entity G port map(lamdaA => P(2)(142),lamdaB => P(2)(398),s => s(2)(142),lamdaOut => P(1)(398));
U_G2399: entity G port map(lamdaA => P(2)(143),lamdaB => P(2)(399),s => s(2)(143),lamdaOut => P(1)(399));
U_G2400: entity G port map(lamdaA => P(2)(144),lamdaB => P(2)(400),s => s(2)(144),lamdaOut => P(1)(400));
U_G2401: entity G port map(lamdaA => P(2)(145),lamdaB => P(2)(401),s => s(2)(145),lamdaOut => P(1)(401));
U_G2402: entity G port map(lamdaA => P(2)(146),lamdaB => P(2)(402),s => s(2)(146),lamdaOut => P(1)(402));
U_G2403: entity G port map(lamdaA => P(2)(147),lamdaB => P(2)(403),s => s(2)(147),lamdaOut => P(1)(403));
U_G2404: entity G port map(lamdaA => P(2)(148),lamdaB => P(2)(404),s => s(2)(148),lamdaOut => P(1)(404));
U_G2405: entity G port map(lamdaA => P(2)(149),lamdaB => P(2)(405),s => s(2)(149),lamdaOut => P(1)(405));
U_G2406: entity G port map(lamdaA => P(2)(150),lamdaB => P(2)(406),s => s(2)(150),lamdaOut => P(1)(406));
U_G2407: entity G port map(lamdaA => P(2)(151),lamdaB => P(2)(407),s => s(2)(151),lamdaOut => P(1)(407));
U_G2408: entity G port map(lamdaA => P(2)(152),lamdaB => P(2)(408),s => s(2)(152),lamdaOut => P(1)(408));
U_G2409: entity G port map(lamdaA => P(2)(153),lamdaB => P(2)(409),s => s(2)(153),lamdaOut => P(1)(409));
U_G2410: entity G port map(lamdaA => P(2)(154),lamdaB => P(2)(410),s => s(2)(154),lamdaOut => P(1)(410));
U_G2411: entity G port map(lamdaA => P(2)(155),lamdaB => P(2)(411),s => s(2)(155),lamdaOut => P(1)(411));
U_G2412: entity G port map(lamdaA => P(2)(156),lamdaB => P(2)(412),s => s(2)(156),lamdaOut => P(1)(412));
U_G2413: entity G port map(lamdaA => P(2)(157),lamdaB => P(2)(413),s => s(2)(157),lamdaOut => P(1)(413));
U_G2414: entity G port map(lamdaA => P(2)(158),lamdaB => P(2)(414),s => s(2)(158),lamdaOut => P(1)(414));
U_G2415: entity G port map(lamdaA => P(2)(159),lamdaB => P(2)(415),s => s(2)(159),lamdaOut => P(1)(415));
U_G2416: entity G port map(lamdaA => P(2)(160),lamdaB => P(2)(416),s => s(2)(160),lamdaOut => P(1)(416));
U_G2417: entity G port map(lamdaA => P(2)(161),lamdaB => P(2)(417),s => s(2)(161),lamdaOut => P(1)(417));
U_G2418: entity G port map(lamdaA => P(2)(162),lamdaB => P(2)(418),s => s(2)(162),lamdaOut => P(1)(418));
U_G2419: entity G port map(lamdaA => P(2)(163),lamdaB => P(2)(419),s => s(2)(163),lamdaOut => P(1)(419));
U_G2420: entity G port map(lamdaA => P(2)(164),lamdaB => P(2)(420),s => s(2)(164),lamdaOut => P(1)(420));
U_G2421: entity G port map(lamdaA => P(2)(165),lamdaB => P(2)(421),s => s(2)(165),lamdaOut => P(1)(421));
U_G2422: entity G port map(lamdaA => P(2)(166),lamdaB => P(2)(422),s => s(2)(166),lamdaOut => P(1)(422));
U_G2423: entity G port map(lamdaA => P(2)(167),lamdaB => P(2)(423),s => s(2)(167),lamdaOut => P(1)(423));
U_G2424: entity G port map(lamdaA => P(2)(168),lamdaB => P(2)(424),s => s(2)(168),lamdaOut => P(1)(424));
U_G2425: entity G port map(lamdaA => P(2)(169),lamdaB => P(2)(425),s => s(2)(169),lamdaOut => P(1)(425));
U_G2426: entity G port map(lamdaA => P(2)(170),lamdaB => P(2)(426),s => s(2)(170),lamdaOut => P(1)(426));
U_G2427: entity G port map(lamdaA => P(2)(171),lamdaB => P(2)(427),s => s(2)(171),lamdaOut => P(1)(427));
U_G2428: entity G port map(lamdaA => P(2)(172),lamdaB => P(2)(428),s => s(2)(172),lamdaOut => P(1)(428));
U_G2429: entity G port map(lamdaA => P(2)(173),lamdaB => P(2)(429),s => s(2)(173),lamdaOut => P(1)(429));
U_G2430: entity G port map(lamdaA => P(2)(174),lamdaB => P(2)(430),s => s(2)(174),lamdaOut => P(1)(430));
U_G2431: entity G port map(lamdaA => P(2)(175),lamdaB => P(2)(431),s => s(2)(175),lamdaOut => P(1)(431));
U_G2432: entity G port map(lamdaA => P(2)(176),lamdaB => P(2)(432),s => s(2)(176),lamdaOut => P(1)(432));
U_G2433: entity G port map(lamdaA => P(2)(177),lamdaB => P(2)(433),s => s(2)(177),lamdaOut => P(1)(433));
U_G2434: entity G port map(lamdaA => P(2)(178),lamdaB => P(2)(434),s => s(2)(178),lamdaOut => P(1)(434));
U_G2435: entity G port map(lamdaA => P(2)(179),lamdaB => P(2)(435),s => s(2)(179),lamdaOut => P(1)(435));
U_G2436: entity G port map(lamdaA => P(2)(180),lamdaB => P(2)(436),s => s(2)(180),lamdaOut => P(1)(436));
U_G2437: entity G port map(lamdaA => P(2)(181),lamdaB => P(2)(437),s => s(2)(181),lamdaOut => P(1)(437));
U_G2438: entity G port map(lamdaA => P(2)(182),lamdaB => P(2)(438),s => s(2)(182),lamdaOut => P(1)(438));
U_G2439: entity G port map(lamdaA => P(2)(183),lamdaB => P(2)(439),s => s(2)(183),lamdaOut => P(1)(439));
U_G2440: entity G port map(lamdaA => P(2)(184),lamdaB => P(2)(440),s => s(2)(184),lamdaOut => P(1)(440));
U_G2441: entity G port map(lamdaA => P(2)(185),lamdaB => P(2)(441),s => s(2)(185),lamdaOut => P(1)(441));
U_G2442: entity G port map(lamdaA => P(2)(186),lamdaB => P(2)(442),s => s(2)(186),lamdaOut => P(1)(442));
U_G2443: entity G port map(lamdaA => P(2)(187),lamdaB => P(2)(443),s => s(2)(187),lamdaOut => P(1)(443));
U_G2444: entity G port map(lamdaA => P(2)(188),lamdaB => P(2)(444),s => s(2)(188),lamdaOut => P(1)(444));
U_G2445: entity G port map(lamdaA => P(2)(189),lamdaB => P(2)(445),s => s(2)(189),lamdaOut => P(1)(445));
U_G2446: entity G port map(lamdaA => P(2)(190),lamdaB => P(2)(446),s => s(2)(190),lamdaOut => P(1)(446));
U_G2447: entity G port map(lamdaA => P(2)(191),lamdaB => P(2)(447),s => s(2)(191),lamdaOut => P(1)(447));
U_G2448: entity G port map(lamdaA => P(2)(192),lamdaB => P(2)(448),s => s(2)(192),lamdaOut => P(1)(448));
U_G2449: entity G port map(lamdaA => P(2)(193),lamdaB => P(2)(449),s => s(2)(193),lamdaOut => P(1)(449));
U_G2450: entity G port map(lamdaA => P(2)(194),lamdaB => P(2)(450),s => s(2)(194),lamdaOut => P(1)(450));
U_G2451: entity G port map(lamdaA => P(2)(195),lamdaB => P(2)(451),s => s(2)(195),lamdaOut => P(1)(451));
U_G2452: entity G port map(lamdaA => P(2)(196),lamdaB => P(2)(452),s => s(2)(196),lamdaOut => P(1)(452));
U_G2453: entity G port map(lamdaA => P(2)(197),lamdaB => P(2)(453),s => s(2)(197),lamdaOut => P(1)(453));
U_G2454: entity G port map(lamdaA => P(2)(198),lamdaB => P(2)(454),s => s(2)(198),lamdaOut => P(1)(454));
U_G2455: entity G port map(lamdaA => P(2)(199),lamdaB => P(2)(455),s => s(2)(199),lamdaOut => P(1)(455));
U_G2456: entity G port map(lamdaA => P(2)(200),lamdaB => P(2)(456),s => s(2)(200),lamdaOut => P(1)(456));
U_G2457: entity G port map(lamdaA => P(2)(201),lamdaB => P(2)(457),s => s(2)(201),lamdaOut => P(1)(457));
U_G2458: entity G port map(lamdaA => P(2)(202),lamdaB => P(2)(458),s => s(2)(202),lamdaOut => P(1)(458));
U_G2459: entity G port map(lamdaA => P(2)(203),lamdaB => P(2)(459),s => s(2)(203),lamdaOut => P(1)(459));
U_G2460: entity G port map(lamdaA => P(2)(204),lamdaB => P(2)(460),s => s(2)(204),lamdaOut => P(1)(460));
U_G2461: entity G port map(lamdaA => P(2)(205),lamdaB => P(2)(461),s => s(2)(205),lamdaOut => P(1)(461));
U_G2462: entity G port map(lamdaA => P(2)(206),lamdaB => P(2)(462),s => s(2)(206),lamdaOut => P(1)(462));
U_G2463: entity G port map(lamdaA => P(2)(207),lamdaB => P(2)(463),s => s(2)(207),lamdaOut => P(1)(463));
U_G2464: entity G port map(lamdaA => P(2)(208),lamdaB => P(2)(464),s => s(2)(208),lamdaOut => P(1)(464));
U_G2465: entity G port map(lamdaA => P(2)(209),lamdaB => P(2)(465),s => s(2)(209),lamdaOut => P(1)(465));
U_G2466: entity G port map(lamdaA => P(2)(210),lamdaB => P(2)(466),s => s(2)(210),lamdaOut => P(1)(466));
U_G2467: entity G port map(lamdaA => P(2)(211),lamdaB => P(2)(467),s => s(2)(211),lamdaOut => P(1)(467));
U_G2468: entity G port map(lamdaA => P(2)(212),lamdaB => P(2)(468),s => s(2)(212),lamdaOut => P(1)(468));
U_G2469: entity G port map(lamdaA => P(2)(213),lamdaB => P(2)(469),s => s(2)(213),lamdaOut => P(1)(469));
U_G2470: entity G port map(lamdaA => P(2)(214),lamdaB => P(2)(470),s => s(2)(214),lamdaOut => P(1)(470));
U_G2471: entity G port map(lamdaA => P(2)(215),lamdaB => P(2)(471),s => s(2)(215),lamdaOut => P(1)(471));
U_G2472: entity G port map(lamdaA => P(2)(216),lamdaB => P(2)(472),s => s(2)(216),lamdaOut => P(1)(472));
U_G2473: entity G port map(lamdaA => P(2)(217),lamdaB => P(2)(473),s => s(2)(217),lamdaOut => P(1)(473));
U_G2474: entity G port map(lamdaA => P(2)(218),lamdaB => P(2)(474),s => s(2)(218),lamdaOut => P(1)(474));
U_G2475: entity G port map(lamdaA => P(2)(219),lamdaB => P(2)(475),s => s(2)(219),lamdaOut => P(1)(475));
U_G2476: entity G port map(lamdaA => P(2)(220),lamdaB => P(2)(476),s => s(2)(220),lamdaOut => P(1)(476));
U_G2477: entity G port map(lamdaA => P(2)(221),lamdaB => P(2)(477),s => s(2)(221),lamdaOut => P(1)(477));
U_G2478: entity G port map(lamdaA => P(2)(222),lamdaB => P(2)(478),s => s(2)(222),lamdaOut => P(1)(478));
U_G2479: entity G port map(lamdaA => P(2)(223),lamdaB => P(2)(479),s => s(2)(223),lamdaOut => P(1)(479));
U_G2480: entity G port map(lamdaA => P(2)(224),lamdaB => P(2)(480),s => s(2)(224),lamdaOut => P(1)(480));
U_G2481: entity G port map(lamdaA => P(2)(225),lamdaB => P(2)(481),s => s(2)(225),lamdaOut => P(1)(481));
U_G2482: entity G port map(lamdaA => P(2)(226),lamdaB => P(2)(482),s => s(2)(226),lamdaOut => P(1)(482));
U_G2483: entity G port map(lamdaA => P(2)(227),lamdaB => P(2)(483),s => s(2)(227),lamdaOut => P(1)(483));
U_G2484: entity G port map(lamdaA => P(2)(228),lamdaB => P(2)(484),s => s(2)(228),lamdaOut => P(1)(484));
U_G2485: entity G port map(lamdaA => P(2)(229),lamdaB => P(2)(485),s => s(2)(229),lamdaOut => P(1)(485));
U_G2486: entity G port map(lamdaA => P(2)(230),lamdaB => P(2)(486),s => s(2)(230),lamdaOut => P(1)(486));
U_G2487: entity G port map(lamdaA => P(2)(231),lamdaB => P(2)(487),s => s(2)(231),lamdaOut => P(1)(487));
U_G2488: entity G port map(lamdaA => P(2)(232),lamdaB => P(2)(488),s => s(2)(232),lamdaOut => P(1)(488));
U_G2489: entity G port map(lamdaA => P(2)(233),lamdaB => P(2)(489),s => s(2)(233),lamdaOut => P(1)(489));
U_G2490: entity G port map(lamdaA => P(2)(234),lamdaB => P(2)(490),s => s(2)(234),lamdaOut => P(1)(490));
U_G2491: entity G port map(lamdaA => P(2)(235),lamdaB => P(2)(491),s => s(2)(235),lamdaOut => P(1)(491));
U_G2492: entity G port map(lamdaA => P(2)(236),lamdaB => P(2)(492),s => s(2)(236),lamdaOut => P(1)(492));
U_G2493: entity G port map(lamdaA => P(2)(237),lamdaB => P(2)(493),s => s(2)(237),lamdaOut => P(1)(493));
U_G2494: entity G port map(lamdaA => P(2)(238),lamdaB => P(2)(494),s => s(2)(238),lamdaOut => P(1)(494));
U_G2495: entity G port map(lamdaA => P(2)(239),lamdaB => P(2)(495),s => s(2)(239),lamdaOut => P(1)(495));
U_G2496: entity G port map(lamdaA => P(2)(240),lamdaB => P(2)(496),s => s(2)(240),lamdaOut => P(1)(496));
U_G2497: entity G port map(lamdaA => P(2)(241),lamdaB => P(2)(497),s => s(2)(241),lamdaOut => P(1)(497));
U_G2498: entity G port map(lamdaA => P(2)(242),lamdaB => P(2)(498),s => s(2)(242),lamdaOut => P(1)(498));
U_G2499: entity G port map(lamdaA => P(2)(243),lamdaB => P(2)(499),s => s(2)(243),lamdaOut => P(1)(499));
U_G2500: entity G port map(lamdaA => P(2)(244),lamdaB => P(2)(500),s => s(2)(244),lamdaOut => P(1)(500));
U_G2501: entity G port map(lamdaA => P(2)(245),lamdaB => P(2)(501),s => s(2)(245),lamdaOut => P(1)(501));
U_G2502: entity G port map(lamdaA => P(2)(246),lamdaB => P(2)(502),s => s(2)(246),lamdaOut => P(1)(502));
U_G2503: entity G port map(lamdaA => P(2)(247),lamdaB => P(2)(503),s => s(2)(247),lamdaOut => P(1)(503));
U_G2504: entity G port map(lamdaA => P(2)(248),lamdaB => P(2)(504),s => s(2)(248),lamdaOut => P(1)(504));
U_G2505: entity G port map(lamdaA => P(2)(249),lamdaB => P(2)(505),s => s(2)(249),lamdaOut => P(1)(505));
U_G2506: entity G port map(lamdaA => P(2)(250),lamdaB => P(2)(506),s => s(2)(250),lamdaOut => P(1)(506));
U_G2507: entity G port map(lamdaA => P(2)(251),lamdaB => P(2)(507),s => s(2)(251),lamdaOut => P(1)(507));
U_G2508: entity G port map(lamdaA => P(2)(252),lamdaB => P(2)(508),s => s(2)(252),lamdaOut => P(1)(508));
U_G2509: entity G port map(lamdaA => P(2)(253),lamdaB => P(2)(509),s => s(2)(253),lamdaOut => P(1)(509));
U_G2510: entity G port map(lamdaA => P(2)(254),lamdaB => P(2)(510),s => s(2)(254),lamdaOut => P(1)(510));
U_G2511: entity G port map(lamdaA => P(2)(255),lamdaB => P(2)(511),s => s(2)(255),lamdaOut => P(1)(511));
U_F2512: entity F port map(lamdaA => P(2)(512),lamdaB => P(2)(768),lamdaOut => P(1)(512));
U_F2513: entity F port map(lamdaA => P(2)(513),lamdaB => P(2)(769),lamdaOut => P(1)(513));
U_F2514: entity F port map(lamdaA => P(2)(514),lamdaB => P(2)(770),lamdaOut => P(1)(514));
U_F2515: entity F port map(lamdaA => P(2)(515),lamdaB => P(2)(771),lamdaOut => P(1)(515));
U_F2516: entity F port map(lamdaA => P(2)(516),lamdaB => P(2)(772),lamdaOut => P(1)(516));
U_F2517: entity F port map(lamdaA => P(2)(517),lamdaB => P(2)(773),lamdaOut => P(1)(517));
U_F2518: entity F port map(lamdaA => P(2)(518),lamdaB => P(2)(774),lamdaOut => P(1)(518));
U_F2519: entity F port map(lamdaA => P(2)(519),lamdaB => P(2)(775),lamdaOut => P(1)(519));
U_F2520: entity F port map(lamdaA => P(2)(520),lamdaB => P(2)(776),lamdaOut => P(1)(520));
U_F2521: entity F port map(lamdaA => P(2)(521),lamdaB => P(2)(777),lamdaOut => P(1)(521));
U_F2522: entity F port map(lamdaA => P(2)(522),lamdaB => P(2)(778),lamdaOut => P(1)(522));
U_F2523: entity F port map(lamdaA => P(2)(523),lamdaB => P(2)(779),lamdaOut => P(1)(523));
U_F2524: entity F port map(lamdaA => P(2)(524),lamdaB => P(2)(780),lamdaOut => P(1)(524));
U_F2525: entity F port map(lamdaA => P(2)(525),lamdaB => P(2)(781),lamdaOut => P(1)(525));
U_F2526: entity F port map(lamdaA => P(2)(526),lamdaB => P(2)(782),lamdaOut => P(1)(526));
U_F2527: entity F port map(lamdaA => P(2)(527),lamdaB => P(2)(783),lamdaOut => P(1)(527));
U_F2528: entity F port map(lamdaA => P(2)(528),lamdaB => P(2)(784),lamdaOut => P(1)(528));
U_F2529: entity F port map(lamdaA => P(2)(529),lamdaB => P(2)(785),lamdaOut => P(1)(529));
U_F2530: entity F port map(lamdaA => P(2)(530),lamdaB => P(2)(786),lamdaOut => P(1)(530));
U_F2531: entity F port map(lamdaA => P(2)(531),lamdaB => P(2)(787),lamdaOut => P(1)(531));
U_F2532: entity F port map(lamdaA => P(2)(532),lamdaB => P(2)(788),lamdaOut => P(1)(532));
U_F2533: entity F port map(lamdaA => P(2)(533),lamdaB => P(2)(789),lamdaOut => P(1)(533));
U_F2534: entity F port map(lamdaA => P(2)(534),lamdaB => P(2)(790),lamdaOut => P(1)(534));
U_F2535: entity F port map(lamdaA => P(2)(535),lamdaB => P(2)(791),lamdaOut => P(1)(535));
U_F2536: entity F port map(lamdaA => P(2)(536),lamdaB => P(2)(792),lamdaOut => P(1)(536));
U_F2537: entity F port map(lamdaA => P(2)(537),lamdaB => P(2)(793),lamdaOut => P(1)(537));
U_F2538: entity F port map(lamdaA => P(2)(538),lamdaB => P(2)(794),lamdaOut => P(1)(538));
U_F2539: entity F port map(lamdaA => P(2)(539),lamdaB => P(2)(795),lamdaOut => P(1)(539));
U_F2540: entity F port map(lamdaA => P(2)(540),lamdaB => P(2)(796),lamdaOut => P(1)(540));
U_F2541: entity F port map(lamdaA => P(2)(541),lamdaB => P(2)(797),lamdaOut => P(1)(541));
U_F2542: entity F port map(lamdaA => P(2)(542),lamdaB => P(2)(798),lamdaOut => P(1)(542));
U_F2543: entity F port map(lamdaA => P(2)(543),lamdaB => P(2)(799),lamdaOut => P(1)(543));
U_F2544: entity F port map(lamdaA => P(2)(544),lamdaB => P(2)(800),lamdaOut => P(1)(544));
U_F2545: entity F port map(lamdaA => P(2)(545),lamdaB => P(2)(801),lamdaOut => P(1)(545));
U_F2546: entity F port map(lamdaA => P(2)(546),lamdaB => P(2)(802),lamdaOut => P(1)(546));
U_F2547: entity F port map(lamdaA => P(2)(547),lamdaB => P(2)(803),lamdaOut => P(1)(547));
U_F2548: entity F port map(lamdaA => P(2)(548),lamdaB => P(2)(804),lamdaOut => P(1)(548));
U_F2549: entity F port map(lamdaA => P(2)(549),lamdaB => P(2)(805),lamdaOut => P(1)(549));
U_F2550: entity F port map(lamdaA => P(2)(550),lamdaB => P(2)(806),lamdaOut => P(1)(550));
U_F2551: entity F port map(lamdaA => P(2)(551),lamdaB => P(2)(807),lamdaOut => P(1)(551));
U_F2552: entity F port map(lamdaA => P(2)(552),lamdaB => P(2)(808),lamdaOut => P(1)(552));
U_F2553: entity F port map(lamdaA => P(2)(553),lamdaB => P(2)(809),lamdaOut => P(1)(553));
U_F2554: entity F port map(lamdaA => P(2)(554),lamdaB => P(2)(810),lamdaOut => P(1)(554));
U_F2555: entity F port map(lamdaA => P(2)(555),lamdaB => P(2)(811),lamdaOut => P(1)(555));
U_F2556: entity F port map(lamdaA => P(2)(556),lamdaB => P(2)(812),lamdaOut => P(1)(556));
U_F2557: entity F port map(lamdaA => P(2)(557),lamdaB => P(2)(813),lamdaOut => P(1)(557));
U_F2558: entity F port map(lamdaA => P(2)(558),lamdaB => P(2)(814),lamdaOut => P(1)(558));
U_F2559: entity F port map(lamdaA => P(2)(559),lamdaB => P(2)(815),lamdaOut => P(1)(559));
U_F2560: entity F port map(lamdaA => P(2)(560),lamdaB => P(2)(816),lamdaOut => P(1)(560));
U_F2561: entity F port map(lamdaA => P(2)(561),lamdaB => P(2)(817),lamdaOut => P(1)(561));
U_F2562: entity F port map(lamdaA => P(2)(562),lamdaB => P(2)(818),lamdaOut => P(1)(562));
U_F2563: entity F port map(lamdaA => P(2)(563),lamdaB => P(2)(819),lamdaOut => P(1)(563));
U_F2564: entity F port map(lamdaA => P(2)(564),lamdaB => P(2)(820),lamdaOut => P(1)(564));
U_F2565: entity F port map(lamdaA => P(2)(565),lamdaB => P(2)(821),lamdaOut => P(1)(565));
U_F2566: entity F port map(lamdaA => P(2)(566),lamdaB => P(2)(822),lamdaOut => P(1)(566));
U_F2567: entity F port map(lamdaA => P(2)(567),lamdaB => P(2)(823),lamdaOut => P(1)(567));
U_F2568: entity F port map(lamdaA => P(2)(568),lamdaB => P(2)(824),lamdaOut => P(1)(568));
U_F2569: entity F port map(lamdaA => P(2)(569),lamdaB => P(2)(825),lamdaOut => P(1)(569));
U_F2570: entity F port map(lamdaA => P(2)(570),lamdaB => P(2)(826),lamdaOut => P(1)(570));
U_F2571: entity F port map(lamdaA => P(2)(571),lamdaB => P(2)(827),lamdaOut => P(1)(571));
U_F2572: entity F port map(lamdaA => P(2)(572),lamdaB => P(2)(828),lamdaOut => P(1)(572));
U_F2573: entity F port map(lamdaA => P(2)(573),lamdaB => P(2)(829),lamdaOut => P(1)(573));
U_F2574: entity F port map(lamdaA => P(2)(574),lamdaB => P(2)(830),lamdaOut => P(1)(574));
U_F2575: entity F port map(lamdaA => P(2)(575),lamdaB => P(2)(831),lamdaOut => P(1)(575));
U_F2576: entity F port map(lamdaA => P(2)(576),lamdaB => P(2)(832),lamdaOut => P(1)(576));
U_F2577: entity F port map(lamdaA => P(2)(577),lamdaB => P(2)(833),lamdaOut => P(1)(577));
U_F2578: entity F port map(lamdaA => P(2)(578),lamdaB => P(2)(834),lamdaOut => P(1)(578));
U_F2579: entity F port map(lamdaA => P(2)(579),lamdaB => P(2)(835),lamdaOut => P(1)(579));
U_F2580: entity F port map(lamdaA => P(2)(580),lamdaB => P(2)(836),lamdaOut => P(1)(580));
U_F2581: entity F port map(lamdaA => P(2)(581),lamdaB => P(2)(837),lamdaOut => P(1)(581));
U_F2582: entity F port map(lamdaA => P(2)(582),lamdaB => P(2)(838),lamdaOut => P(1)(582));
U_F2583: entity F port map(lamdaA => P(2)(583),lamdaB => P(2)(839),lamdaOut => P(1)(583));
U_F2584: entity F port map(lamdaA => P(2)(584),lamdaB => P(2)(840),lamdaOut => P(1)(584));
U_F2585: entity F port map(lamdaA => P(2)(585),lamdaB => P(2)(841),lamdaOut => P(1)(585));
U_F2586: entity F port map(lamdaA => P(2)(586),lamdaB => P(2)(842),lamdaOut => P(1)(586));
U_F2587: entity F port map(lamdaA => P(2)(587),lamdaB => P(2)(843),lamdaOut => P(1)(587));
U_F2588: entity F port map(lamdaA => P(2)(588),lamdaB => P(2)(844),lamdaOut => P(1)(588));
U_F2589: entity F port map(lamdaA => P(2)(589),lamdaB => P(2)(845),lamdaOut => P(1)(589));
U_F2590: entity F port map(lamdaA => P(2)(590),lamdaB => P(2)(846),lamdaOut => P(1)(590));
U_F2591: entity F port map(lamdaA => P(2)(591),lamdaB => P(2)(847),lamdaOut => P(1)(591));
U_F2592: entity F port map(lamdaA => P(2)(592),lamdaB => P(2)(848),lamdaOut => P(1)(592));
U_F2593: entity F port map(lamdaA => P(2)(593),lamdaB => P(2)(849),lamdaOut => P(1)(593));
U_F2594: entity F port map(lamdaA => P(2)(594),lamdaB => P(2)(850),lamdaOut => P(1)(594));
U_F2595: entity F port map(lamdaA => P(2)(595),lamdaB => P(2)(851),lamdaOut => P(1)(595));
U_F2596: entity F port map(lamdaA => P(2)(596),lamdaB => P(2)(852),lamdaOut => P(1)(596));
U_F2597: entity F port map(lamdaA => P(2)(597),lamdaB => P(2)(853),lamdaOut => P(1)(597));
U_F2598: entity F port map(lamdaA => P(2)(598),lamdaB => P(2)(854),lamdaOut => P(1)(598));
U_F2599: entity F port map(lamdaA => P(2)(599),lamdaB => P(2)(855),lamdaOut => P(1)(599));
U_F2600: entity F port map(lamdaA => P(2)(600),lamdaB => P(2)(856),lamdaOut => P(1)(600));
U_F2601: entity F port map(lamdaA => P(2)(601),lamdaB => P(2)(857),lamdaOut => P(1)(601));
U_F2602: entity F port map(lamdaA => P(2)(602),lamdaB => P(2)(858),lamdaOut => P(1)(602));
U_F2603: entity F port map(lamdaA => P(2)(603),lamdaB => P(2)(859),lamdaOut => P(1)(603));
U_F2604: entity F port map(lamdaA => P(2)(604),lamdaB => P(2)(860),lamdaOut => P(1)(604));
U_F2605: entity F port map(lamdaA => P(2)(605),lamdaB => P(2)(861),lamdaOut => P(1)(605));
U_F2606: entity F port map(lamdaA => P(2)(606),lamdaB => P(2)(862),lamdaOut => P(1)(606));
U_F2607: entity F port map(lamdaA => P(2)(607),lamdaB => P(2)(863),lamdaOut => P(1)(607));
U_F2608: entity F port map(lamdaA => P(2)(608),lamdaB => P(2)(864),lamdaOut => P(1)(608));
U_F2609: entity F port map(lamdaA => P(2)(609),lamdaB => P(2)(865),lamdaOut => P(1)(609));
U_F2610: entity F port map(lamdaA => P(2)(610),lamdaB => P(2)(866),lamdaOut => P(1)(610));
U_F2611: entity F port map(lamdaA => P(2)(611),lamdaB => P(2)(867),lamdaOut => P(1)(611));
U_F2612: entity F port map(lamdaA => P(2)(612),lamdaB => P(2)(868),lamdaOut => P(1)(612));
U_F2613: entity F port map(lamdaA => P(2)(613),lamdaB => P(2)(869),lamdaOut => P(1)(613));
U_F2614: entity F port map(lamdaA => P(2)(614),lamdaB => P(2)(870),lamdaOut => P(1)(614));
U_F2615: entity F port map(lamdaA => P(2)(615),lamdaB => P(2)(871),lamdaOut => P(1)(615));
U_F2616: entity F port map(lamdaA => P(2)(616),lamdaB => P(2)(872),lamdaOut => P(1)(616));
U_F2617: entity F port map(lamdaA => P(2)(617),lamdaB => P(2)(873),lamdaOut => P(1)(617));
U_F2618: entity F port map(lamdaA => P(2)(618),lamdaB => P(2)(874),lamdaOut => P(1)(618));
U_F2619: entity F port map(lamdaA => P(2)(619),lamdaB => P(2)(875),lamdaOut => P(1)(619));
U_F2620: entity F port map(lamdaA => P(2)(620),lamdaB => P(2)(876),lamdaOut => P(1)(620));
U_F2621: entity F port map(lamdaA => P(2)(621),lamdaB => P(2)(877),lamdaOut => P(1)(621));
U_F2622: entity F port map(lamdaA => P(2)(622),lamdaB => P(2)(878),lamdaOut => P(1)(622));
U_F2623: entity F port map(lamdaA => P(2)(623),lamdaB => P(2)(879),lamdaOut => P(1)(623));
U_F2624: entity F port map(lamdaA => P(2)(624),lamdaB => P(2)(880),lamdaOut => P(1)(624));
U_F2625: entity F port map(lamdaA => P(2)(625),lamdaB => P(2)(881),lamdaOut => P(1)(625));
U_F2626: entity F port map(lamdaA => P(2)(626),lamdaB => P(2)(882),lamdaOut => P(1)(626));
U_F2627: entity F port map(lamdaA => P(2)(627),lamdaB => P(2)(883),lamdaOut => P(1)(627));
U_F2628: entity F port map(lamdaA => P(2)(628),lamdaB => P(2)(884),lamdaOut => P(1)(628));
U_F2629: entity F port map(lamdaA => P(2)(629),lamdaB => P(2)(885),lamdaOut => P(1)(629));
U_F2630: entity F port map(lamdaA => P(2)(630),lamdaB => P(2)(886),lamdaOut => P(1)(630));
U_F2631: entity F port map(lamdaA => P(2)(631),lamdaB => P(2)(887),lamdaOut => P(1)(631));
U_F2632: entity F port map(lamdaA => P(2)(632),lamdaB => P(2)(888),lamdaOut => P(1)(632));
U_F2633: entity F port map(lamdaA => P(2)(633),lamdaB => P(2)(889),lamdaOut => P(1)(633));
U_F2634: entity F port map(lamdaA => P(2)(634),lamdaB => P(2)(890),lamdaOut => P(1)(634));
U_F2635: entity F port map(lamdaA => P(2)(635),lamdaB => P(2)(891),lamdaOut => P(1)(635));
U_F2636: entity F port map(lamdaA => P(2)(636),lamdaB => P(2)(892),lamdaOut => P(1)(636));
U_F2637: entity F port map(lamdaA => P(2)(637),lamdaB => P(2)(893),lamdaOut => P(1)(637));
U_F2638: entity F port map(lamdaA => P(2)(638),lamdaB => P(2)(894),lamdaOut => P(1)(638));
U_F2639: entity F port map(lamdaA => P(2)(639),lamdaB => P(2)(895),lamdaOut => P(1)(639));
U_F2640: entity F port map(lamdaA => P(2)(640),lamdaB => P(2)(896),lamdaOut => P(1)(640));
U_F2641: entity F port map(lamdaA => P(2)(641),lamdaB => P(2)(897),lamdaOut => P(1)(641));
U_F2642: entity F port map(lamdaA => P(2)(642),lamdaB => P(2)(898),lamdaOut => P(1)(642));
U_F2643: entity F port map(lamdaA => P(2)(643),lamdaB => P(2)(899),lamdaOut => P(1)(643));
U_F2644: entity F port map(lamdaA => P(2)(644),lamdaB => P(2)(900),lamdaOut => P(1)(644));
U_F2645: entity F port map(lamdaA => P(2)(645),lamdaB => P(2)(901),lamdaOut => P(1)(645));
U_F2646: entity F port map(lamdaA => P(2)(646),lamdaB => P(2)(902),lamdaOut => P(1)(646));
U_F2647: entity F port map(lamdaA => P(2)(647),lamdaB => P(2)(903),lamdaOut => P(1)(647));
U_F2648: entity F port map(lamdaA => P(2)(648),lamdaB => P(2)(904),lamdaOut => P(1)(648));
U_F2649: entity F port map(lamdaA => P(2)(649),lamdaB => P(2)(905),lamdaOut => P(1)(649));
U_F2650: entity F port map(lamdaA => P(2)(650),lamdaB => P(2)(906),lamdaOut => P(1)(650));
U_F2651: entity F port map(lamdaA => P(2)(651),lamdaB => P(2)(907),lamdaOut => P(1)(651));
U_F2652: entity F port map(lamdaA => P(2)(652),lamdaB => P(2)(908),lamdaOut => P(1)(652));
U_F2653: entity F port map(lamdaA => P(2)(653),lamdaB => P(2)(909),lamdaOut => P(1)(653));
U_F2654: entity F port map(lamdaA => P(2)(654),lamdaB => P(2)(910),lamdaOut => P(1)(654));
U_F2655: entity F port map(lamdaA => P(2)(655),lamdaB => P(2)(911),lamdaOut => P(1)(655));
U_F2656: entity F port map(lamdaA => P(2)(656),lamdaB => P(2)(912),lamdaOut => P(1)(656));
U_F2657: entity F port map(lamdaA => P(2)(657),lamdaB => P(2)(913),lamdaOut => P(1)(657));
U_F2658: entity F port map(lamdaA => P(2)(658),lamdaB => P(2)(914),lamdaOut => P(1)(658));
U_F2659: entity F port map(lamdaA => P(2)(659),lamdaB => P(2)(915),lamdaOut => P(1)(659));
U_F2660: entity F port map(lamdaA => P(2)(660),lamdaB => P(2)(916),lamdaOut => P(1)(660));
U_F2661: entity F port map(lamdaA => P(2)(661),lamdaB => P(2)(917),lamdaOut => P(1)(661));
U_F2662: entity F port map(lamdaA => P(2)(662),lamdaB => P(2)(918),lamdaOut => P(1)(662));
U_F2663: entity F port map(lamdaA => P(2)(663),lamdaB => P(2)(919),lamdaOut => P(1)(663));
U_F2664: entity F port map(lamdaA => P(2)(664),lamdaB => P(2)(920),lamdaOut => P(1)(664));
U_F2665: entity F port map(lamdaA => P(2)(665),lamdaB => P(2)(921),lamdaOut => P(1)(665));
U_F2666: entity F port map(lamdaA => P(2)(666),lamdaB => P(2)(922),lamdaOut => P(1)(666));
U_F2667: entity F port map(lamdaA => P(2)(667),lamdaB => P(2)(923),lamdaOut => P(1)(667));
U_F2668: entity F port map(lamdaA => P(2)(668),lamdaB => P(2)(924),lamdaOut => P(1)(668));
U_F2669: entity F port map(lamdaA => P(2)(669),lamdaB => P(2)(925),lamdaOut => P(1)(669));
U_F2670: entity F port map(lamdaA => P(2)(670),lamdaB => P(2)(926),lamdaOut => P(1)(670));
U_F2671: entity F port map(lamdaA => P(2)(671),lamdaB => P(2)(927),lamdaOut => P(1)(671));
U_F2672: entity F port map(lamdaA => P(2)(672),lamdaB => P(2)(928),lamdaOut => P(1)(672));
U_F2673: entity F port map(lamdaA => P(2)(673),lamdaB => P(2)(929),lamdaOut => P(1)(673));
U_F2674: entity F port map(lamdaA => P(2)(674),lamdaB => P(2)(930),lamdaOut => P(1)(674));
U_F2675: entity F port map(lamdaA => P(2)(675),lamdaB => P(2)(931),lamdaOut => P(1)(675));
U_F2676: entity F port map(lamdaA => P(2)(676),lamdaB => P(2)(932),lamdaOut => P(1)(676));
U_F2677: entity F port map(lamdaA => P(2)(677),lamdaB => P(2)(933),lamdaOut => P(1)(677));
U_F2678: entity F port map(lamdaA => P(2)(678),lamdaB => P(2)(934),lamdaOut => P(1)(678));
U_F2679: entity F port map(lamdaA => P(2)(679),lamdaB => P(2)(935),lamdaOut => P(1)(679));
U_F2680: entity F port map(lamdaA => P(2)(680),lamdaB => P(2)(936),lamdaOut => P(1)(680));
U_F2681: entity F port map(lamdaA => P(2)(681),lamdaB => P(2)(937),lamdaOut => P(1)(681));
U_F2682: entity F port map(lamdaA => P(2)(682),lamdaB => P(2)(938),lamdaOut => P(1)(682));
U_F2683: entity F port map(lamdaA => P(2)(683),lamdaB => P(2)(939),lamdaOut => P(1)(683));
U_F2684: entity F port map(lamdaA => P(2)(684),lamdaB => P(2)(940),lamdaOut => P(1)(684));
U_F2685: entity F port map(lamdaA => P(2)(685),lamdaB => P(2)(941),lamdaOut => P(1)(685));
U_F2686: entity F port map(lamdaA => P(2)(686),lamdaB => P(2)(942),lamdaOut => P(1)(686));
U_F2687: entity F port map(lamdaA => P(2)(687),lamdaB => P(2)(943),lamdaOut => P(1)(687));
U_F2688: entity F port map(lamdaA => P(2)(688),lamdaB => P(2)(944),lamdaOut => P(1)(688));
U_F2689: entity F port map(lamdaA => P(2)(689),lamdaB => P(2)(945),lamdaOut => P(1)(689));
U_F2690: entity F port map(lamdaA => P(2)(690),lamdaB => P(2)(946),lamdaOut => P(1)(690));
U_F2691: entity F port map(lamdaA => P(2)(691),lamdaB => P(2)(947),lamdaOut => P(1)(691));
U_F2692: entity F port map(lamdaA => P(2)(692),lamdaB => P(2)(948),lamdaOut => P(1)(692));
U_F2693: entity F port map(lamdaA => P(2)(693),lamdaB => P(2)(949),lamdaOut => P(1)(693));
U_F2694: entity F port map(lamdaA => P(2)(694),lamdaB => P(2)(950),lamdaOut => P(1)(694));
U_F2695: entity F port map(lamdaA => P(2)(695),lamdaB => P(2)(951),lamdaOut => P(1)(695));
U_F2696: entity F port map(lamdaA => P(2)(696),lamdaB => P(2)(952),lamdaOut => P(1)(696));
U_F2697: entity F port map(lamdaA => P(2)(697),lamdaB => P(2)(953),lamdaOut => P(1)(697));
U_F2698: entity F port map(lamdaA => P(2)(698),lamdaB => P(2)(954),lamdaOut => P(1)(698));
U_F2699: entity F port map(lamdaA => P(2)(699),lamdaB => P(2)(955),lamdaOut => P(1)(699));
U_F2700: entity F port map(lamdaA => P(2)(700),lamdaB => P(2)(956),lamdaOut => P(1)(700));
U_F2701: entity F port map(lamdaA => P(2)(701),lamdaB => P(2)(957),lamdaOut => P(1)(701));
U_F2702: entity F port map(lamdaA => P(2)(702),lamdaB => P(2)(958),lamdaOut => P(1)(702));
U_F2703: entity F port map(lamdaA => P(2)(703),lamdaB => P(2)(959),lamdaOut => P(1)(703));
U_F2704: entity F port map(lamdaA => P(2)(704),lamdaB => P(2)(960),lamdaOut => P(1)(704));
U_F2705: entity F port map(lamdaA => P(2)(705),lamdaB => P(2)(961),lamdaOut => P(1)(705));
U_F2706: entity F port map(lamdaA => P(2)(706),lamdaB => P(2)(962),lamdaOut => P(1)(706));
U_F2707: entity F port map(lamdaA => P(2)(707),lamdaB => P(2)(963),lamdaOut => P(1)(707));
U_F2708: entity F port map(lamdaA => P(2)(708),lamdaB => P(2)(964),lamdaOut => P(1)(708));
U_F2709: entity F port map(lamdaA => P(2)(709),lamdaB => P(2)(965),lamdaOut => P(1)(709));
U_F2710: entity F port map(lamdaA => P(2)(710),lamdaB => P(2)(966),lamdaOut => P(1)(710));
U_F2711: entity F port map(lamdaA => P(2)(711),lamdaB => P(2)(967),lamdaOut => P(1)(711));
U_F2712: entity F port map(lamdaA => P(2)(712),lamdaB => P(2)(968),lamdaOut => P(1)(712));
U_F2713: entity F port map(lamdaA => P(2)(713),lamdaB => P(2)(969),lamdaOut => P(1)(713));
U_F2714: entity F port map(lamdaA => P(2)(714),lamdaB => P(2)(970),lamdaOut => P(1)(714));
U_F2715: entity F port map(lamdaA => P(2)(715),lamdaB => P(2)(971),lamdaOut => P(1)(715));
U_F2716: entity F port map(lamdaA => P(2)(716),lamdaB => P(2)(972),lamdaOut => P(1)(716));
U_F2717: entity F port map(lamdaA => P(2)(717),lamdaB => P(2)(973),lamdaOut => P(1)(717));
U_F2718: entity F port map(lamdaA => P(2)(718),lamdaB => P(2)(974),lamdaOut => P(1)(718));
U_F2719: entity F port map(lamdaA => P(2)(719),lamdaB => P(2)(975),lamdaOut => P(1)(719));
U_F2720: entity F port map(lamdaA => P(2)(720),lamdaB => P(2)(976),lamdaOut => P(1)(720));
U_F2721: entity F port map(lamdaA => P(2)(721),lamdaB => P(2)(977),lamdaOut => P(1)(721));
U_F2722: entity F port map(lamdaA => P(2)(722),lamdaB => P(2)(978),lamdaOut => P(1)(722));
U_F2723: entity F port map(lamdaA => P(2)(723),lamdaB => P(2)(979),lamdaOut => P(1)(723));
U_F2724: entity F port map(lamdaA => P(2)(724),lamdaB => P(2)(980),lamdaOut => P(1)(724));
U_F2725: entity F port map(lamdaA => P(2)(725),lamdaB => P(2)(981),lamdaOut => P(1)(725));
U_F2726: entity F port map(lamdaA => P(2)(726),lamdaB => P(2)(982),lamdaOut => P(1)(726));
U_F2727: entity F port map(lamdaA => P(2)(727),lamdaB => P(2)(983),lamdaOut => P(1)(727));
U_F2728: entity F port map(lamdaA => P(2)(728),lamdaB => P(2)(984),lamdaOut => P(1)(728));
U_F2729: entity F port map(lamdaA => P(2)(729),lamdaB => P(2)(985),lamdaOut => P(1)(729));
U_F2730: entity F port map(lamdaA => P(2)(730),lamdaB => P(2)(986),lamdaOut => P(1)(730));
U_F2731: entity F port map(lamdaA => P(2)(731),lamdaB => P(2)(987),lamdaOut => P(1)(731));
U_F2732: entity F port map(lamdaA => P(2)(732),lamdaB => P(2)(988),lamdaOut => P(1)(732));
U_F2733: entity F port map(lamdaA => P(2)(733),lamdaB => P(2)(989),lamdaOut => P(1)(733));
U_F2734: entity F port map(lamdaA => P(2)(734),lamdaB => P(2)(990),lamdaOut => P(1)(734));
U_F2735: entity F port map(lamdaA => P(2)(735),lamdaB => P(2)(991),lamdaOut => P(1)(735));
U_F2736: entity F port map(lamdaA => P(2)(736),lamdaB => P(2)(992),lamdaOut => P(1)(736));
U_F2737: entity F port map(lamdaA => P(2)(737),lamdaB => P(2)(993),lamdaOut => P(1)(737));
U_F2738: entity F port map(lamdaA => P(2)(738),lamdaB => P(2)(994),lamdaOut => P(1)(738));
U_F2739: entity F port map(lamdaA => P(2)(739),lamdaB => P(2)(995),lamdaOut => P(1)(739));
U_F2740: entity F port map(lamdaA => P(2)(740),lamdaB => P(2)(996),lamdaOut => P(1)(740));
U_F2741: entity F port map(lamdaA => P(2)(741),lamdaB => P(2)(997),lamdaOut => P(1)(741));
U_F2742: entity F port map(lamdaA => P(2)(742),lamdaB => P(2)(998),lamdaOut => P(1)(742));
U_F2743: entity F port map(lamdaA => P(2)(743),lamdaB => P(2)(999),lamdaOut => P(1)(743));
U_F2744: entity F port map(lamdaA => P(2)(744),lamdaB => P(2)(1000),lamdaOut => P(1)(744));
U_F2745: entity F port map(lamdaA => P(2)(745),lamdaB => P(2)(1001),lamdaOut => P(1)(745));
U_F2746: entity F port map(lamdaA => P(2)(746),lamdaB => P(2)(1002),lamdaOut => P(1)(746));
U_F2747: entity F port map(lamdaA => P(2)(747),lamdaB => P(2)(1003),lamdaOut => P(1)(747));
U_F2748: entity F port map(lamdaA => P(2)(748),lamdaB => P(2)(1004),lamdaOut => P(1)(748));
U_F2749: entity F port map(lamdaA => P(2)(749),lamdaB => P(2)(1005),lamdaOut => P(1)(749));
U_F2750: entity F port map(lamdaA => P(2)(750),lamdaB => P(2)(1006),lamdaOut => P(1)(750));
U_F2751: entity F port map(lamdaA => P(2)(751),lamdaB => P(2)(1007),lamdaOut => P(1)(751));
U_F2752: entity F port map(lamdaA => P(2)(752),lamdaB => P(2)(1008),lamdaOut => P(1)(752));
U_F2753: entity F port map(lamdaA => P(2)(753),lamdaB => P(2)(1009),lamdaOut => P(1)(753));
U_F2754: entity F port map(lamdaA => P(2)(754),lamdaB => P(2)(1010),lamdaOut => P(1)(754));
U_F2755: entity F port map(lamdaA => P(2)(755),lamdaB => P(2)(1011),lamdaOut => P(1)(755));
U_F2756: entity F port map(lamdaA => P(2)(756),lamdaB => P(2)(1012),lamdaOut => P(1)(756));
U_F2757: entity F port map(lamdaA => P(2)(757),lamdaB => P(2)(1013),lamdaOut => P(1)(757));
U_F2758: entity F port map(lamdaA => P(2)(758),lamdaB => P(2)(1014),lamdaOut => P(1)(758));
U_F2759: entity F port map(lamdaA => P(2)(759),lamdaB => P(2)(1015),lamdaOut => P(1)(759));
U_F2760: entity F port map(lamdaA => P(2)(760),lamdaB => P(2)(1016),lamdaOut => P(1)(760));
U_F2761: entity F port map(lamdaA => P(2)(761),lamdaB => P(2)(1017),lamdaOut => P(1)(761));
U_F2762: entity F port map(lamdaA => P(2)(762),lamdaB => P(2)(1018),lamdaOut => P(1)(762));
U_F2763: entity F port map(lamdaA => P(2)(763),lamdaB => P(2)(1019),lamdaOut => P(1)(763));
U_F2764: entity F port map(lamdaA => P(2)(764),lamdaB => P(2)(1020),lamdaOut => P(1)(764));
U_F2765: entity F port map(lamdaA => P(2)(765),lamdaB => P(2)(1021),lamdaOut => P(1)(765));
U_F2766: entity F port map(lamdaA => P(2)(766),lamdaB => P(2)(1022),lamdaOut => P(1)(766));
U_F2767: entity F port map(lamdaA => P(2)(767),lamdaB => P(2)(1023),lamdaOut => P(1)(767));
U_G2768: entity G port map(lamdaA => P(2)(512),lamdaB => P(2)(768),s => s(2)(256),lamdaOut => P(1)(768));
U_G2769: entity G port map(lamdaA => P(2)(513),lamdaB => P(2)(769),s => s(2)(257),lamdaOut => P(1)(769));
U_G2770: entity G port map(lamdaA => P(2)(514),lamdaB => P(2)(770),s => s(2)(258),lamdaOut => P(1)(770));
U_G2771: entity G port map(lamdaA => P(2)(515),lamdaB => P(2)(771),s => s(2)(259),lamdaOut => P(1)(771));
U_G2772: entity G port map(lamdaA => P(2)(516),lamdaB => P(2)(772),s => s(2)(260),lamdaOut => P(1)(772));
U_G2773: entity G port map(lamdaA => P(2)(517),lamdaB => P(2)(773),s => s(2)(261),lamdaOut => P(1)(773));
U_G2774: entity G port map(lamdaA => P(2)(518),lamdaB => P(2)(774),s => s(2)(262),lamdaOut => P(1)(774));
U_G2775: entity G port map(lamdaA => P(2)(519),lamdaB => P(2)(775),s => s(2)(263),lamdaOut => P(1)(775));
U_G2776: entity G port map(lamdaA => P(2)(520),lamdaB => P(2)(776),s => s(2)(264),lamdaOut => P(1)(776));
U_G2777: entity G port map(lamdaA => P(2)(521),lamdaB => P(2)(777),s => s(2)(265),lamdaOut => P(1)(777));
U_G2778: entity G port map(lamdaA => P(2)(522),lamdaB => P(2)(778),s => s(2)(266),lamdaOut => P(1)(778));
U_G2779: entity G port map(lamdaA => P(2)(523),lamdaB => P(2)(779),s => s(2)(267),lamdaOut => P(1)(779));
U_G2780: entity G port map(lamdaA => P(2)(524),lamdaB => P(2)(780),s => s(2)(268),lamdaOut => P(1)(780));
U_G2781: entity G port map(lamdaA => P(2)(525),lamdaB => P(2)(781),s => s(2)(269),lamdaOut => P(1)(781));
U_G2782: entity G port map(lamdaA => P(2)(526),lamdaB => P(2)(782),s => s(2)(270),lamdaOut => P(1)(782));
U_G2783: entity G port map(lamdaA => P(2)(527),lamdaB => P(2)(783),s => s(2)(271),lamdaOut => P(1)(783));
U_G2784: entity G port map(lamdaA => P(2)(528),lamdaB => P(2)(784),s => s(2)(272),lamdaOut => P(1)(784));
U_G2785: entity G port map(lamdaA => P(2)(529),lamdaB => P(2)(785),s => s(2)(273),lamdaOut => P(1)(785));
U_G2786: entity G port map(lamdaA => P(2)(530),lamdaB => P(2)(786),s => s(2)(274),lamdaOut => P(1)(786));
U_G2787: entity G port map(lamdaA => P(2)(531),lamdaB => P(2)(787),s => s(2)(275),lamdaOut => P(1)(787));
U_G2788: entity G port map(lamdaA => P(2)(532),lamdaB => P(2)(788),s => s(2)(276),lamdaOut => P(1)(788));
U_G2789: entity G port map(lamdaA => P(2)(533),lamdaB => P(2)(789),s => s(2)(277),lamdaOut => P(1)(789));
U_G2790: entity G port map(lamdaA => P(2)(534),lamdaB => P(2)(790),s => s(2)(278),lamdaOut => P(1)(790));
U_G2791: entity G port map(lamdaA => P(2)(535),lamdaB => P(2)(791),s => s(2)(279),lamdaOut => P(1)(791));
U_G2792: entity G port map(lamdaA => P(2)(536),lamdaB => P(2)(792),s => s(2)(280),lamdaOut => P(1)(792));
U_G2793: entity G port map(lamdaA => P(2)(537),lamdaB => P(2)(793),s => s(2)(281),lamdaOut => P(1)(793));
U_G2794: entity G port map(lamdaA => P(2)(538),lamdaB => P(2)(794),s => s(2)(282),lamdaOut => P(1)(794));
U_G2795: entity G port map(lamdaA => P(2)(539),lamdaB => P(2)(795),s => s(2)(283),lamdaOut => P(1)(795));
U_G2796: entity G port map(lamdaA => P(2)(540),lamdaB => P(2)(796),s => s(2)(284),lamdaOut => P(1)(796));
U_G2797: entity G port map(lamdaA => P(2)(541),lamdaB => P(2)(797),s => s(2)(285),lamdaOut => P(1)(797));
U_G2798: entity G port map(lamdaA => P(2)(542),lamdaB => P(2)(798),s => s(2)(286),lamdaOut => P(1)(798));
U_G2799: entity G port map(lamdaA => P(2)(543),lamdaB => P(2)(799),s => s(2)(287),lamdaOut => P(1)(799));
U_G2800: entity G port map(lamdaA => P(2)(544),lamdaB => P(2)(800),s => s(2)(288),lamdaOut => P(1)(800));
U_G2801: entity G port map(lamdaA => P(2)(545),lamdaB => P(2)(801),s => s(2)(289),lamdaOut => P(1)(801));
U_G2802: entity G port map(lamdaA => P(2)(546),lamdaB => P(2)(802),s => s(2)(290),lamdaOut => P(1)(802));
U_G2803: entity G port map(lamdaA => P(2)(547),lamdaB => P(2)(803),s => s(2)(291),lamdaOut => P(1)(803));
U_G2804: entity G port map(lamdaA => P(2)(548),lamdaB => P(2)(804),s => s(2)(292),lamdaOut => P(1)(804));
U_G2805: entity G port map(lamdaA => P(2)(549),lamdaB => P(2)(805),s => s(2)(293),lamdaOut => P(1)(805));
U_G2806: entity G port map(lamdaA => P(2)(550),lamdaB => P(2)(806),s => s(2)(294),lamdaOut => P(1)(806));
U_G2807: entity G port map(lamdaA => P(2)(551),lamdaB => P(2)(807),s => s(2)(295),lamdaOut => P(1)(807));
U_G2808: entity G port map(lamdaA => P(2)(552),lamdaB => P(2)(808),s => s(2)(296),lamdaOut => P(1)(808));
U_G2809: entity G port map(lamdaA => P(2)(553),lamdaB => P(2)(809),s => s(2)(297),lamdaOut => P(1)(809));
U_G2810: entity G port map(lamdaA => P(2)(554),lamdaB => P(2)(810),s => s(2)(298),lamdaOut => P(1)(810));
U_G2811: entity G port map(lamdaA => P(2)(555),lamdaB => P(2)(811),s => s(2)(299),lamdaOut => P(1)(811));
U_G2812: entity G port map(lamdaA => P(2)(556),lamdaB => P(2)(812),s => s(2)(300),lamdaOut => P(1)(812));
U_G2813: entity G port map(lamdaA => P(2)(557),lamdaB => P(2)(813),s => s(2)(301),lamdaOut => P(1)(813));
U_G2814: entity G port map(lamdaA => P(2)(558),lamdaB => P(2)(814),s => s(2)(302),lamdaOut => P(1)(814));
U_G2815: entity G port map(lamdaA => P(2)(559),lamdaB => P(2)(815),s => s(2)(303),lamdaOut => P(1)(815));
U_G2816: entity G port map(lamdaA => P(2)(560),lamdaB => P(2)(816),s => s(2)(304),lamdaOut => P(1)(816));
U_G2817: entity G port map(lamdaA => P(2)(561),lamdaB => P(2)(817),s => s(2)(305),lamdaOut => P(1)(817));
U_G2818: entity G port map(lamdaA => P(2)(562),lamdaB => P(2)(818),s => s(2)(306),lamdaOut => P(1)(818));
U_G2819: entity G port map(lamdaA => P(2)(563),lamdaB => P(2)(819),s => s(2)(307),lamdaOut => P(1)(819));
U_G2820: entity G port map(lamdaA => P(2)(564),lamdaB => P(2)(820),s => s(2)(308),lamdaOut => P(1)(820));
U_G2821: entity G port map(lamdaA => P(2)(565),lamdaB => P(2)(821),s => s(2)(309),lamdaOut => P(1)(821));
U_G2822: entity G port map(lamdaA => P(2)(566),lamdaB => P(2)(822),s => s(2)(310),lamdaOut => P(1)(822));
U_G2823: entity G port map(lamdaA => P(2)(567),lamdaB => P(2)(823),s => s(2)(311),lamdaOut => P(1)(823));
U_G2824: entity G port map(lamdaA => P(2)(568),lamdaB => P(2)(824),s => s(2)(312),lamdaOut => P(1)(824));
U_G2825: entity G port map(lamdaA => P(2)(569),lamdaB => P(2)(825),s => s(2)(313),lamdaOut => P(1)(825));
U_G2826: entity G port map(lamdaA => P(2)(570),lamdaB => P(2)(826),s => s(2)(314),lamdaOut => P(1)(826));
U_G2827: entity G port map(lamdaA => P(2)(571),lamdaB => P(2)(827),s => s(2)(315),lamdaOut => P(1)(827));
U_G2828: entity G port map(lamdaA => P(2)(572),lamdaB => P(2)(828),s => s(2)(316),lamdaOut => P(1)(828));
U_G2829: entity G port map(lamdaA => P(2)(573),lamdaB => P(2)(829),s => s(2)(317),lamdaOut => P(1)(829));
U_G2830: entity G port map(lamdaA => P(2)(574),lamdaB => P(2)(830),s => s(2)(318),lamdaOut => P(1)(830));
U_G2831: entity G port map(lamdaA => P(2)(575),lamdaB => P(2)(831),s => s(2)(319),lamdaOut => P(1)(831));
U_G2832: entity G port map(lamdaA => P(2)(576),lamdaB => P(2)(832),s => s(2)(320),lamdaOut => P(1)(832));
U_G2833: entity G port map(lamdaA => P(2)(577),lamdaB => P(2)(833),s => s(2)(321),lamdaOut => P(1)(833));
U_G2834: entity G port map(lamdaA => P(2)(578),lamdaB => P(2)(834),s => s(2)(322),lamdaOut => P(1)(834));
U_G2835: entity G port map(lamdaA => P(2)(579),lamdaB => P(2)(835),s => s(2)(323),lamdaOut => P(1)(835));
U_G2836: entity G port map(lamdaA => P(2)(580),lamdaB => P(2)(836),s => s(2)(324),lamdaOut => P(1)(836));
U_G2837: entity G port map(lamdaA => P(2)(581),lamdaB => P(2)(837),s => s(2)(325),lamdaOut => P(1)(837));
U_G2838: entity G port map(lamdaA => P(2)(582),lamdaB => P(2)(838),s => s(2)(326),lamdaOut => P(1)(838));
U_G2839: entity G port map(lamdaA => P(2)(583),lamdaB => P(2)(839),s => s(2)(327),lamdaOut => P(1)(839));
U_G2840: entity G port map(lamdaA => P(2)(584),lamdaB => P(2)(840),s => s(2)(328),lamdaOut => P(1)(840));
U_G2841: entity G port map(lamdaA => P(2)(585),lamdaB => P(2)(841),s => s(2)(329),lamdaOut => P(1)(841));
U_G2842: entity G port map(lamdaA => P(2)(586),lamdaB => P(2)(842),s => s(2)(330),lamdaOut => P(1)(842));
U_G2843: entity G port map(lamdaA => P(2)(587),lamdaB => P(2)(843),s => s(2)(331),lamdaOut => P(1)(843));
U_G2844: entity G port map(lamdaA => P(2)(588),lamdaB => P(2)(844),s => s(2)(332),lamdaOut => P(1)(844));
U_G2845: entity G port map(lamdaA => P(2)(589),lamdaB => P(2)(845),s => s(2)(333),lamdaOut => P(1)(845));
U_G2846: entity G port map(lamdaA => P(2)(590),lamdaB => P(2)(846),s => s(2)(334),lamdaOut => P(1)(846));
U_G2847: entity G port map(lamdaA => P(2)(591),lamdaB => P(2)(847),s => s(2)(335),lamdaOut => P(1)(847));
U_G2848: entity G port map(lamdaA => P(2)(592),lamdaB => P(2)(848),s => s(2)(336),lamdaOut => P(1)(848));
U_G2849: entity G port map(lamdaA => P(2)(593),lamdaB => P(2)(849),s => s(2)(337),lamdaOut => P(1)(849));
U_G2850: entity G port map(lamdaA => P(2)(594),lamdaB => P(2)(850),s => s(2)(338),lamdaOut => P(1)(850));
U_G2851: entity G port map(lamdaA => P(2)(595),lamdaB => P(2)(851),s => s(2)(339),lamdaOut => P(1)(851));
U_G2852: entity G port map(lamdaA => P(2)(596),lamdaB => P(2)(852),s => s(2)(340),lamdaOut => P(1)(852));
U_G2853: entity G port map(lamdaA => P(2)(597),lamdaB => P(2)(853),s => s(2)(341),lamdaOut => P(1)(853));
U_G2854: entity G port map(lamdaA => P(2)(598),lamdaB => P(2)(854),s => s(2)(342),lamdaOut => P(1)(854));
U_G2855: entity G port map(lamdaA => P(2)(599),lamdaB => P(2)(855),s => s(2)(343),lamdaOut => P(1)(855));
U_G2856: entity G port map(lamdaA => P(2)(600),lamdaB => P(2)(856),s => s(2)(344),lamdaOut => P(1)(856));
U_G2857: entity G port map(lamdaA => P(2)(601),lamdaB => P(2)(857),s => s(2)(345),lamdaOut => P(1)(857));
U_G2858: entity G port map(lamdaA => P(2)(602),lamdaB => P(2)(858),s => s(2)(346),lamdaOut => P(1)(858));
U_G2859: entity G port map(lamdaA => P(2)(603),lamdaB => P(2)(859),s => s(2)(347),lamdaOut => P(1)(859));
U_G2860: entity G port map(lamdaA => P(2)(604),lamdaB => P(2)(860),s => s(2)(348),lamdaOut => P(1)(860));
U_G2861: entity G port map(lamdaA => P(2)(605),lamdaB => P(2)(861),s => s(2)(349),lamdaOut => P(1)(861));
U_G2862: entity G port map(lamdaA => P(2)(606),lamdaB => P(2)(862),s => s(2)(350),lamdaOut => P(1)(862));
U_G2863: entity G port map(lamdaA => P(2)(607),lamdaB => P(2)(863),s => s(2)(351),lamdaOut => P(1)(863));
U_G2864: entity G port map(lamdaA => P(2)(608),lamdaB => P(2)(864),s => s(2)(352),lamdaOut => P(1)(864));
U_G2865: entity G port map(lamdaA => P(2)(609),lamdaB => P(2)(865),s => s(2)(353),lamdaOut => P(1)(865));
U_G2866: entity G port map(lamdaA => P(2)(610),lamdaB => P(2)(866),s => s(2)(354),lamdaOut => P(1)(866));
U_G2867: entity G port map(lamdaA => P(2)(611),lamdaB => P(2)(867),s => s(2)(355),lamdaOut => P(1)(867));
U_G2868: entity G port map(lamdaA => P(2)(612),lamdaB => P(2)(868),s => s(2)(356),lamdaOut => P(1)(868));
U_G2869: entity G port map(lamdaA => P(2)(613),lamdaB => P(2)(869),s => s(2)(357),lamdaOut => P(1)(869));
U_G2870: entity G port map(lamdaA => P(2)(614),lamdaB => P(2)(870),s => s(2)(358),lamdaOut => P(1)(870));
U_G2871: entity G port map(lamdaA => P(2)(615),lamdaB => P(2)(871),s => s(2)(359),lamdaOut => P(1)(871));
U_G2872: entity G port map(lamdaA => P(2)(616),lamdaB => P(2)(872),s => s(2)(360),lamdaOut => P(1)(872));
U_G2873: entity G port map(lamdaA => P(2)(617),lamdaB => P(2)(873),s => s(2)(361),lamdaOut => P(1)(873));
U_G2874: entity G port map(lamdaA => P(2)(618),lamdaB => P(2)(874),s => s(2)(362),lamdaOut => P(1)(874));
U_G2875: entity G port map(lamdaA => P(2)(619),lamdaB => P(2)(875),s => s(2)(363),lamdaOut => P(1)(875));
U_G2876: entity G port map(lamdaA => P(2)(620),lamdaB => P(2)(876),s => s(2)(364),lamdaOut => P(1)(876));
U_G2877: entity G port map(lamdaA => P(2)(621),lamdaB => P(2)(877),s => s(2)(365),lamdaOut => P(1)(877));
U_G2878: entity G port map(lamdaA => P(2)(622),lamdaB => P(2)(878),s => s(2)(366),lamdaOut => P(1)(878));
U_G2879: entity G port map(lamdaA => P(2)(623),lamdaB => P(2)(879),s => s(2)(367),lamdaOut => P(1)(879));
U_G2880: entity G port map(lamdaA => P(2)(624),lamdaB => P(2)(880),s => s(2)(368),lamdaOut => P(1)(880));
U_G2881: entity G port map(lamdaA => P(2)(625),lamdaB => P(2)(881),s => s(2)(369),lamdaOut => P(1)(881));
U_G2882: entity G port map(lamdaA => P(2)(626),lamdaB => P(2)(882),s => s(2)(370),lamdaOut => P(1)(882));
U_G2883: entity G port map(lamdaA => P(2)(627),lamdaB => P(2)(883),s => s(2)(371),lamdaOut => P(1)(883));
U_G2884: entity G port map(lamdaA => P(2)(628),lamdaB => P(2)(884),s => s(2)(372),lamdaOut => P(1)(884));
U_G2885: entity G port map(lamdaA => P(2)(629),lamdaB => P(2)(885),s => s(2)(373),lamdaOut => P(1)(885));
U_G2886: entity G port map(lamdaA => P(2)(630),lamdaB => P(2)(886),s => s(2)(374),lamdaOut => P(1)(886));
U_G2887: entity G port map(lamdaA => P(2)(631),lamdaB => P(2)(887),s => s(2)(375),lamdaOut => P(1)(887));
U_G2888: entity G port map(lamdaA => P(2)(632),lamdaB => P(2)(888),s => s(2)(376),lamdaOut => P(1)(888));
U_G2889: entity G port map(lamdaA => P(2)(633),lamdaB => P(2)(889),s => s(2)(377),lamdaOut => P(1)(889));
U_G2890: entity G port map(lamdaA => P(2)(634),lamdaB => P(2)(890),s => s(2)(378),lamdaOut => P(1)(890));
U_G2891: entity G port map(lamdaA => P(2)(635),lamdaB => P(2)(891),s => s(2)(379),lamdaOut => P(1)(891));
U_G2892: entity G port map(lamdaA => P(2)(636),lamdaB => P(2)(892),s => s(2)(380),lamdaOut => P(1)(892));
U_G2893: entity G port map(lamdaA => P(2)(637),lamdaB => P(2)(893),s => s(2)(381),lamdaOut => P(1)(893));
U_G2894: entity G port map(lamdaA => P(2)(638),lamdaB => P(2)(894),s => s(2)(382),lamdaOut => P(1)(894));
U_G2895: entity G port map(lamdaA => P(2)(639),lamdaB => P(2)(895),s => s(2)(383),lamdaOut => P(1)(895));
U_G2896: entity G port map(lamdaA => P(2)(640),lamdaB => P(2)(896),s => s(2)(384),lamdaOut => P(1)(896));
U_G2897: entity G port map(lamdaA => P(2)(641),lamdaB => P(2)(897),s => s(2)(385),lamdaOut => P(1)(897));
U_G2898: entity G port map(lamdaA => P(2)(642),lamdaB => P(2)(898),s => s(2)(386),lamdaOut => P(1)(898));
U_G2899: entity G port map(lamdaA => P(2)(643),lamdaB => P(2)(899),s => s(2)(387),lamdaOut => P(1)(899));
U_G2900: entity G port map(lamdaA => P(2)(644),lamdaB => P(2)(900),s => s(2)(388),lamdaOut => P(1)(900));
U_G2901: entity G port map(lamdaA => P(2)(645),lamdaB => P(2)(901),s => s(2)(389),lamdaOut => P(1)(901));
U_G2902: entity G port map(lamdaA => P(2)(646),lamdaB => P(2)(902),s => s(2)(390),lamdaOut => P(1)(902));
U_G2903: entity G port map(lamdaA => P(2)(647),lamdaB => P(2)(903),s => s(2)(391),lamdaOut => P(1)(903));
U_G2904: entity G port map(lamdaA => P(2)(648),lamdaB => P(2)(904),s => s(2)(392),lamdaOut => P(1)(904));
U_G2905: entity G port map(lamdaA => P(2)(649),lamdaB => P(2)(905),s => s(2)(393),lamdaOut => P(1)(905));
U_G2906: entity G port map(lamdaA => P(2)(650),lamdaB => P(2)(906),s => s(2)(394),lamdaOut => P(1)(906));
U_G2907: entity G port map(lamdaA => P(2)(651),lamdaB => P(2)(907),s => s(2)(395),lamdaOut => P(1)(907));
U_G2908: entity G port map(lamdaA => P(2)(652),lamdaB => P(2)(908),s => s(2)(396),lamdaOut => P(1)(908));
U_G2909: entity G port map(lamdaA => P(2)(653),lamdaB => P(2)(909),s => s(2)(397),lamdaOut => P(1)(909));
U_G2910: entity G port map(lamdaA => P(2)(654),lamdaB => P(2)(910),s => s(2)(398),lamdaOut => P(1)(910));
U_G2911: entity G port map(lamdaA => P(2)(655),lamdaB => P(2)(911),s => s(2)(399),lamdaOut => P(1)(911));
U_G2912: entity G port map(lamdaA => P(2)(656),lamdaB => P(2)(912),s => s(2)(400),lamdaOut => P(1)(912));
U_G2913: entity G port map(lamdaA => P(2)(657),lamdaB => P(2)(913),s => s(2)(401),lamdaOut => P(1)(913));
U_G2914: entity G port map(lamdaA => P(2)(658),lamdaB => P(2)(914),s => s(2)(402),lamdaOut => P(1)(914));
U_G2915: entity G port map(lamdaA => P(2)(659),lamdaB => P(2)(915),s => s(2)(403),lamdaOut => P(1)(915));
U_G2916: entity G port map(lamdaA => P(2)(660),lamdaB => P(2)(916),s => s(2)(404),lamdaOut => P(1)(916));
U_G2917: entity G port map(lamdaA => P(2)(661),lamdaB => P(2)(917),s => s(2)(405),lamdaOut => P(1)(917));
U_G2918: entity G port map(lamdaA => P(2)(662),lamdaB => P(2)(918),s => s(2)(406),lamdaOut => P(1)(918));
U_G2919: entity G port map(lamdaA => P(2)(663),lamdaB => P(2)(919),s => s(2)(407),lamdaOut => P(1)(919));
U_G2920: entity G port map(lamdaA => P(2)(664),lamdaB => P(2)(920),s => s(2)(408),lamdaOut => P(1)(920));
U_G2921: entity G port map(lamdaA => P(2)(665),lamdaB => P(2)(921),s => s(2)(409),lamdaOut => P(1)(921));
U_G2922: entity G port map(lamdaA => P(2)(666),lamdaB => P(2)(922),s => s(2)(410),lamdaOut => P(1)(922));
U_G2923: entity G port map(lamdaA => P(2)(667),lamdaB => P(2)(923),s => s(2)(411),lamdaOut => P(1)(923));
U_G2924: entity G port map(lamdaA => P(2)(668),lamdaB => P(2)(924),s => s(2)(412),lamdaOut => P(1)(924));
U_G2925: entity G port map(lamdaA => P(2)(669),lamdaB => P(2)(925),s => s(2)(413),lamdaOut => P(1)(925));
U_G2926: entity G port map(lamdaA => P(2)(670),lamdaB => P(2)(926),s => s(2)(414),lamdaOut => P(1)(926));
U_G2927: entity G port map(lamdaA => P(2)(671),lamdaB => P(2)(927),s => s(2)(415),lamdaOut => P(1)(927));
U_G2928: entity G port map(lamdaA => P(2)(672),lamdaB => P(2)(928),s => s(2)(416),lamdaOut => P(1)(928));
U_G2929: entity G port map(lamdaA => P(2)(673),lamdaB => P(2)(929),s => s(2)(417),lamdaOut => P(1)(929));
U_G2930: entity G port map(lamdaA => P(2)(674),lamdaB => P(2)(930),s => s(2)(418),lamdaOut => P(1)(930));
U_G2931: entity G port map(lamdaA => P(2)(675),lamdaB => P(2)(931),s => s(2)(419),lamdaOut => P(1)(931));
U_G2932: entity G port map(lamdaA => P(2)(676),lamdaB => P(2)(932),s => s(2)(420),lamdaOut => P(1)(932));
U_G2933: entity G port map(lamdaA => P(2)(677),lamdaB => P(2)(933),s => s(2)(421),lamdaOut => P(1)(933));
U_G2934: entity G port map(lamdaA => P(2)(678),lamdaB => P(2)(934),s => s(2)(422),lamdaOut => P(1)(934));
U_G2935: entity G port map(lamdaA => P(2)(679),lamdaB => P(2)(935),s => s(2)(423),lamdaOut => P(1)(935));
U_G2936: entity G port map(lamdaA => P(2)(680),lamdaB => P(2)(936),s => s(2)(424),lamdaOut => P(1)(936));
U_G2937: entity G port map(lamdaA => P(2)(681),lamdaB => P(2)(937),s => s(2)(425),lamdaOut => P(1)(937));
U_G2938: entity G port map(lamdaA => P(2)(682),lamdaB => P(2)(938),s => s(2)(426),lamdaOut => P(1)(938));
U_G2939: entity G port map(lamdaA => P(2)(683),lamdaB => P(2)(939),s => s(2)(427),lamdaOut => P(1)(939));
U_G2940: entity G port map(lamdaA => P(2)(684),lamdaB => P(2)(940),s => s(2)(428),lamdaOut => P(1)(940));
U_G2941: entity G port map(lamdaA => P(2)(685),lamdaB => P(2)(941),s => s(2)(429),lamdaOut => P(1)(941));
U_G2942: entity G port map(lamdaA => P(2)(686),lamdaB => P(2)(942),s => s(2)(430),lamdaOut => P(1)(942));
U_G2943: entity G port map(lamdaA => P(2)(687),lamdaB => P(2)(943),s => s(2)(431),lamdaOut => P(1)(943));
U_G2944: entity G port map(lamdaA => P(2)(688),lamdaB => P(2)(944),s => s(2)(432),lamdaOut => P(1)(944));
U_G2945: entity G port map(lamdaA => P(2)(689),lamdaB => P(2)(945),s => s(2)(433),lamdaOut => P(1)(945));
U_G2946: entity G port map(lamdaA => P(2)(690),lamdaB => P(2)(946),s => s(2)(434),lamdaOut => P(1)(946));
U_G2947: entity G port map(lamdaA => P(2)(691),lamdaB => P(2)(947),s => s(2)(435),lamdaOut => P(1)(947));
U_G2948: entity G port map(lamdaA => P(2)(692),lamdaB => P(2)(948),s => s(2)(436),lamdaOut => P(1)(948));
U_G2949: entity G port map(lamdaA => P(2)(693),lamdaB => P(2)(949),s => s(2)(437),lamdaOut => P(1)(949));
U_G2950: entity G port map(lamdaA => P(2)(694),lamdaB => P(2)(950),s => s(2)(438),lamdaOut => P(1)(950));
U_G2951: entity G port map(lamdaA => P(2)(695),lamdaB => P(2)(951),s => s(2)(439),lamdaOut => P(1)(951));
U_G2952: entity G port map(lamdaA => P(2)(696),lamdaB => P(2)(952),s => s(2)(440),lamdaOut => P(1)(952));
U_G2953: entity G port map(lamdaA => P(2)(697),lamdaB => P(2)(953),s => s(2)(441),lamdaOut => P(1)(953));
U_G2954: entity G port map(lamdaA => P(2)(698),lamdaB => P(2)(954),s => s(2)(442),lamdaOut => P(1)(954));
U_G2955: entity G port map(lamdaA => P(2)(699),lamdaB => P(2)(955),s => s(2)(443),lamdaOut => P(1)(955));
U_G2956: entity G port map(lamdaA => P(2)(700),lamdaB => P(2)(956),s => s(2)(444),lamdaOut => P(1)(956));
U_G2957: entity G port map(lamdaA => P(2)(701),lamdaB => P(2)(957),s => s(2)(445),lamdaOut => P(1)(957));
U_G2958: entity G port map(lamdaA => P(2)(702),lamdaB => P(2)(958),s => s(2)(446),lamdaOut => P(1)(958));
U_G2959: entity G port map(lamdaA => P(2)(703),lamdaB => P(2)(959),s => s(2)(447),lamdaOut => P(1)(959));
U_G2960: entity G port map(lamdaA => P(2)(704),lamdaB => P(2)(960),s => s(2)(448),lamdaOut => P(1)(960));
U_G2961: entity G port map(lamdaA => P(2)(705),lamdaB => P(2)(961),s => s(2)(449),lamdaOut => P(1)(961));
U_G2962: entity G port map(lamdaA => P(2)(706),lamdaB => P(2)(962),s => s(2)(450),lamdaOut => P(1)(962));
U_G2963: entity G port map(lamdaA => P(2)(707),lamdaB => P(2)(963),s => s(2)(451),lamdaOut => P(1)(963));
U_G2964: entity G port map(lamdaA => P(2)(708),lamdaB => P(2)(964),s => s(2)(452),lamdaOut => P(1)(964));
U_G2965: entity G port map(lamdaA => P(2)(709),lamdaB => P(2)(965),s => s(2)(453),lamdaOut => P(1)(965));
U_G2966: entity G port map(lamdaA => P(2)(710),lamdaB => P(2)(966),s => s(2)(454),lamdaOut => P(1)(966));
U_G2967: entity G port map(lamdaA => P(2)(711),lamdaB => P(2)(967),s => s(2)(455),lamdaOut => P(1)(967));
U_G2968: entity G port map(lamdaA => P(2)(712),lamdaB => P(2)(968),s => s(2)(456),lamdaOut => P(1)(968));
U_G2969: entity G port map(lamdaA => P(2)(713),lamdaB => P(2)(969),s => s(2)(457),lamdaOut => P(1)(969));
U_G2970: entity G port map(lamdaA => P(2)(714),lamdaB => P(2)(970),s => s(2)(458),lamdaOut => P(1)(970));
U_G2971: entity G port map(lamdaA => P(2)(715),lamdaB => P(2)(971),s => s(2)(459),lamdaOut => P(1)(971));
U_G2972: entity G port map(lamdaA => P(2)(716),lamdaB => P(2)(972),s => s(2)(460),lamdaOut => P(1)(972));
U_G2973: entity G port map(lamdaA => P(2)(717),lamdaB => P(2)(973),s => s(2)(461),lamdaOut => P(1)(973));
U_G2974: entity G port map(lamdaA => P(2)(718),lamdaB => P(2)(974),s => s(2)(462),lamdaOut => P(1)(974));
U_G2975: entity G port map(lamdaA => P(2)(719),lamdaB => P(2)(975),s => s(2)(463),lamdaOut => P(1)(975));
U_G2976: entity G port map(lamdaA => P(2)(720),lamdaB => P(2)(976),s => s(2)(464),lamdaOut => P(1)(976));
U_G2977: entity G port map(lamdaA => P(2)(721),lamdaB => P(2)(977),s => s(2)(465),lamdaOut => P(1)(977));
U_G2978: entity G port map(lamdaA => P(2)(722),lamdaB => P(2)(978),s => s(2)(466),lamdaOut => P(1)(978));
U_G2979: entity G port map(lamdaA => P(2)(723),lamdaB => P(2)(979),s => s(2)(467),lamdaOut => P(1)(979));
U_G2980: entity G port map(lamdaA => P(2)(724),lamdaB => P(2)(980),s => s(2)(468),lamdaOut => P(1)(980));
U_G2981: entity G port map(lamdaA => P(2)(725),lamdaB => P(2)(981),s => s(2)(469),lamdaOut => P(1)(981));
U_G2982: entity G port map(lamdaA => P(2)(726),lamdaB => P(2)(982),s => s(2)(470),lamdaOut => P(1)(982));
U_G2983: entity G port map(lamdaA => P(2)(727),lamdaB => P(2)(983),s => s(2)(471),lamdaOut => P(1)(983));
U_G2984: entity G port map(lamdaA => P(2)(728),lamdaB => P(2)(984),s => s(2)(472),lamdaOut => P(1)(984));
U_G2985: entity G port map(lamdaA => P(2)(729),lamdaB => P(2)(985),s => s(2)(473),lamdaOut => P(1)(985));
U_G2986: entity G port map(lamdaA => P(2)(730),lamdaB => P(2)(986),s => s(2)(474),lamdaOut => P(1)(986));
U_G2987: entity G port map(lamdaA => P(2)(731),lamdaB => P(2)(987),s => s(2)(475),lamdaOut => P(1)(987));
U_G2988: entity G port map(lamdaA => P(2)(732),lamdaB => P(2)(988),s => s(2)(476),lamdaOut => P(1)(988));
U_G2989: entity G port map(lamdaA => P(2)(733),lamdaB => P(2)(989),s => s(2)(477),lamdaOut => P(1)(989));
U_G2990: entity G port map(lamdaA => P(2)(734),lamdaB => P(2)(990),s => s(2)(478),lamdaOut => P(1)(990));
U_G2991: entity G port map(lamdaA => P(2)(735),lamdaB => P(2)(991),s => s(2)(479),lamdaOut => P(1)(991));
U_G2992: entity G port map(lamdaA => P(2)(736),lamdaB => P(2)(992),s => s(2)(480),lamdaOut => P(1)(992));
U_G2993: entity G port map(lamdaA => P(2)(737),lamdaB => P(2)(993),s => s(2)(481),lamdaOut => P(1)(993));
U_G2994: entity G port map(lamdaA => P(2)(738),lamdaB => P(2)(994),s => s(2)(482),lamdaOut => P(1)(994));
U_G2995: entity G port map(lamdaA => P(2)(739),lamdaB => P(2)(995),s => s(2)(483),lamdaOut => P(1)(995));
U_G2996: entity G port map(lamdaA => P(2)(740),lamdaB => P(2)(996),s => s(2)(484),lamdaOut => P(1)(996));
U_G2997: entity G port map(lamdaA => P(2)(741),lamdaB => P(2)(997),s => s(2)(485),lamdaOut => P(1)(997));
U_G2998: entity G port map(lamdaA => P(2)(742),lamdaB => P(2)(998),s => s(2)(486),lamdaOut => P(1)(998));
U_G2999: entity G port map(lamdaA => P(2)(743),lamdaB => P(2)(999),s => s(2)(487),lamdaOut => P(1)(999));
U_G21000: entity G port map(lamdaA => P(2)(744),lamdaB => P(2)(1000),s => s(2)(488),lamdaOut => P(1)(1000));
U_G21001: entity G port map(lamdaA => P(2)(745),lamdaB => P(2)(1001),s => s(2)(489),lamdaOut => P(1)(1001));
U_G21002: entity G port map(lamdaA => P(2)(746),lamdaB => P(2)(1002),s => s(2)(490),lamdaOut => P(1)(1002));
U_G21003: entity G port map(lamdaA => P(2)(747),lamdaB => P(2)(1003),s => s(2)(491),lamdaOut => P(1)(1003));
U_G21004: entity G port map(lamdaA => P(2)(748),lamdaB => P(2)(1004),s => s(2)(492),lamdaOut => P(1)(1004));
U_G21005: entity G port map(lamdaA => P(2)(749),lamdaB => P(2)(1005),s => s(2)(493),lamdaOut => P(1)(1005));
U_G21006: entity G port map(lamdaA => P(2)(750),lamdaB => P(2)(1006),s => s(2)(494),lamdaOut => P(1)(1006));
U_G21007: entity G port map(lamdaA => P(2)(751),lamdaB => P(2)(1007),s => s(2)(495),lamdaOut => P(1)(1007));
U_G21008: entity G port map(lamdaA => P(2)(752),lamdaB => P(2)(1008),s => s(2)(496),lamdaOut => P(1)(1008));
U_G21009: entity G port map(lamdaA => P(2)(753),lamdaB => P(2)(1009),s => s(2)(497),lamdaOut => P(1)(1009));
U_G21010: entity G port map(lamdaA => P(2)(754),lamdaB => P(2)(1010),s => s(2)(498),lamdaOut => P(1)(1010));
U_G21011: entity G port map(lamdaA => P(2)(755),lamdaB => P(2)(1011),s => s(2)(499),lamdaOut => P(1)(1011));
U_G21012: entity G port map(lamdaA => P(2)(756),lamdaB => P(2)(1012),s => s(2)(500),lamdaOut => P(1)(1012));
U_G21013: entity G port map(lamdaA => P(2)(757),lamdaB => P(2)(1013),s => s(2)(501),lamdaOut => P(1)(1013));
U_G21014: entity G port map(lamdaA => P(2)(758),lamdaB => P(2)(1014),s => s(2)(502),lamdaOut => P(1)(1014));
U_G21015: entity G port map(lamdaA => P(2)(759),lamdaB => P(2)(1015),s => s(2)(503),lamdaOut => P(1)(1015));
U_G21016: entity G port map(lamdaA => P(2)(760),lamdaB => P(2)(1016),s => s(2)(504),lamdaOut => P(1)(1016));
U_G21017: entity G port map(lamdaA => P(2)(761),lamdaB => P(2)(1017),s => s(2)(505),lamdaOut => P(1)(1017));
U_G21018: entity G port map(lamdaA => P(2)(762),lamdaB => P(2)(1018),s => s(2)(506),lamdaOut => P(1)(1018));
U_G21019: entity G port map(lamdaA => P(2)(763),lamdaB => P(2)(1019),s => s(2)(507),lamdaOut => P(1)(1019));
U_G21020: entity G port map(lamdaA => P(2)(764),lamdaB => P(2)(1020),s => s(2)(508),lamdaOut => P(1)(1020));
U_G21021: entity G port map(lamdaA => P(2)(765),lamdaB => P(2)(1021),s => s(2)(509),lamdaOut => P(1)(1021));
U_G21022: entity G port map(lamdaA => P(2)(766),lamdaB => P(2)(1022),s => s(2)(510),lamdaOut => P(1)(1022));
U_G21023: entity G port map(lamdaA => P(2)(767),lamdaB => P(2)(1023),s => s(2)(511),lamdaOut => P(1)(1023));
-- STAGE 0
U_F10: entity F port map(lamdaA => P(1)(0),lamdaB => P(1)(512),lamdaOut => P(0)(0));
U_F11: entity F port map(lamdaA => P(1)(1),lamdaB => P(1)(513),lamdaOut => P(0)(1));
U_F12: entity F port map(lamdaA => P(1)(2),lamdaB => P(1)(514),lamdaOut => P(0)(2));
U_F13: entity F port map(lamdaA => P(1)(3),lamdaB => P(1)(515),lamdaOut => P(0)(3));
U_F14: entity F port map(lamdaA => P(1)(4),lamdaB => P(1)(516),lamdaOut => P(0)(4));
U_F15: entity F port map(lamdaA => P(1)(5),lamdaB => P(1)(517),lamdaOut => P(0)(5));
U_F16: entity F port map(lamdaA => P(1)(6),lamdaB => P(1)(518),lamdaOut => P(0)(6));
U_F17: entity F port map(lamdaA => P(1)(7),lamdaB => P(1)(519),lamdaOut => P(0)(7));
U_F18: entity F port map(lamdaA => P(1)(8),lamdaB => P(1)(520),lamdaOut => P(0)(8));
U_F19: entity F port map(lamdaA => P(1)(9),lamdaB => P(1)(521),lamdaOut => P(0)(9));
U_F110: entity F port map(lamdaA => P(1)(10),lamdaB => P(1)(522),lamdaOut => P(0)(10));
U_F111: entity F port map(lamdaA => P(1)(11),lamdaB => P(1)(523),lamdaOut => P(0)(11));
U_F112: entity F port map(lamdaA => P(1)(12),lamdaB => P(1)(524),lamdaOut => P(0)(12));
U_F113: entity F port map(lamdaA => P(1)(13),lamdaB => P(1)(525),lamdaOut => P(0)(13));
U_F114: entity F port map(lamdaA => P(1)(14),lamdaB => P(1)(526),lamdaOut => P(0)(14));
U_F115: entity F port map(lamdaA => P(1)(15),lamdaB => P(1)(527),lamdaOut => P(0)(15));
U_F116: entity F port map(lamdaA => P(1)(16),lamdaB => P(1)(528),lamdaOut => P(0)(16));
U_F117: entity F port map(lamdaA => P(1)(17),lamdaB => P(1)(529),lamdaOut => P(0)(17));
U_F118: entity F port map(lamdaA => P(1)(18),lamdaB => P(1)(530),lamdaOut => P(0)(18));
U_F119: entity F port map(lamdaA => P(1)(19),lamdaB => P(1)(531),lamdaOut => P(0)(19));
U_F120: entity F port map(lamdaA => P(1)(20),lamdaB => P(1)(532),lamdaOut => P(0)(20));
U_F121: entity F port map(lamdaA => P(1)(21),lamdaB => P(1)(533),lamdaOut => P(0)(21));
U_F122: entity F port map(lamdaA => P(1)(22),lamdaB => P(1)(534),lamdaOut => P(0)(22));
U_F123: entity F port map(lamdaA => P(1)(23),lamdaB => P(1)(535),lamdaOut => P(0)(23));
U_F124: entity F port map(lamdaA => P(1)(24),lamdaB => P(1)(536),lamdaOut => P(0)(24));
U_F125: entity F port map(lamdaA => P(1)(25),lamdaB => P(1)(537),lamdaOut => P(0)(25));
U_F126: entity F port map(lamdaA => P(1)(26),lamdaB => P(1)(538),lamdaOut => P(0)(26));
U_F127: entity F port map(lamdaA => P(1)(27),lamdaB => P(1)(539),lamdaOut => P(0)(27));
U_F128: entity F port map(lamdaA => P(1)(28),lamdaB => P(1)(540),lamdaOut => P(0)(28));
U_F129: entity F port map(lamdaA => P(1)(29),lamdaB => P(1)(541),lamdaOut => P(0)(29));
U_F130: entity F port map(lamdaA => P(1)(30),lamdaB => P(1)(542),lamdaOut => P(0)(30));
U_F131: entity F port map(lamdaA => P(1)(31),lamdaB => P(1)(543),lamdaOut => P(0)(31));
U_F132: entity F port map(lamdaA => P(1)(32),lamdaB => P(1)(544),lamdaOut => P(0)(32));
U_F133: entity F port map(lamdaA => P(1)(33),lamdaB => P(1)(545),lamdaOut => P(0)(33));
U_F134: entity F port map(lamdaA => P(1)(34),lamdaB => P(1)(546),lamdaOut => P(0)(34));
U_F135: entity F port map(lamdaA => P(1)(35),lamdaB => P(1)(547),lamdaOut => P(0)(35));
U_F136: entity F port map(lamdaA => P(1)(36),lamdaB => P(1)(548),lamdaOut => P(0)(36));
U_F137: entity F port map(lamdaA => P(1)(37),lamdaB => P(1)(549),lamdaOut => P(0)(37));
U_F138: entity F port map(lamdaA => P(1)(38),lamdaB => P(1)(550),lamdaOut => P(0)(38));
U_F139: entity F port map(lamdaA => P(1)(39),lamdaB => P(1)(551),lamdaOut => P(0)(39));
U_F140: entity F port map(lamdaA => P(1)(40),lamdaB => P(1)(552),lamdaOut => P(0)(40));
U_F141: entity F port map(lamdaA => P(1)(41),lamdaB => P(1)(553),lamdaOut => P(0)(41));
U_F142: entity F port map(lamdaA => P(1)(42),lamdaB => P(1)(554),lamdaOut => P(0)(42));
U_F143: entity F port map(lamdaA => P(1)(43),lamdaB => P(1)(555),lamdaOut => P(0)(43));
U_F144: entity F port map(lamdaA => P(1)(44),lamdaB => P(1)(556),lamdaOut => P(0)(44));
U_F145: entity F port map(lamdaA => P(1)(45),lamdaB => P(1)(557),lamdaOut => P(0)(45));
U_F146: entity F port map(lamdaA => P(1)(46),lamdaB => P(1)(558),lamdaOut => P(0)(46));
U_F147: entity F port map(lamdaA => P(1)(47),lamdaB => P(1)(559),lamdaOut => P(0)(47));
U_F148: entity F port map(lamdaA => P(1)(48),lamdaB => P(1)(560),lamdaOut => P(0)(48));
U_F149: entity F port map(lamdaA => P(1)(49),lamdaB => P(1)(561),lamdaOut => P(0)(49));
U_F150: entity F port map(lamdaA => P(1)(50),lamdaB => P(1)(562),lamdaOut => P(0)(50));
U_F151: entity F port map(lamdaA => P(1)(51),lamdaB => P(1)(563),lamdaOut => P(0)(51));
U_F152: entity F port map(lamdaA => P(1)(52),lamdaB => P(1)(564),lamdaOut => P(0)(52));
U_F153: entity F port map(lamdaA => P(1)(53),lamdaB => P(1)(565),lamdaOut => P(0)(53));
U_F154: entity F port map(lamdaA => P(1)(54),lamdaB => P(1)(566),lamdaOut => P(0)(54));
U_F155: entity F port map(lamdaA => P(1)(55),lamdaB => P(1)(567),lamdaOut => P(0)(55));
U_F156: entity F port map(lamdaA => P(1)(56),lamdaB => P(1)(568),lamdaOut => P(0)(56));
U_F157: entity F port map(lamdaA => P(1)(57),lamdaB => P(1)(569),lamdaOut => P(0)(57));
U_F158: entity F port map(lamdaA => P(1)(58),lamdaB => P(1)(570),lamdaOut => P(0)(58));
U_F159: entity F port map(lamdaA => P(1)(59),lamdaB => P(1)(571),lamdaOut => P(0)(59));
U_F160: entity F port map(lamdaA => P(1)(60),lamdaB => P(1)(572),lamdaOut => P(0)(60));
U_F161: entity F port map(lamdaA => P(1)(61),lamdaB => P(1)(573),lamdaOut => P(0)(61));
U_F162: entity F port map(lamdaA => P(1)(62),lamdaB => P(1)(574),lamdaOut => P(0)(62));
U_F163: entity F port map(lamdaA => P(1)(63),lamdaB => P(1)(575),lamdaOut => P(0)(63));
U_F164: entity F port map(lamdaA => P(1)(64),lamdaB => P(1)(576),lamdaOut => P(0)(64));
U_F165: entity F port map(lamdaA => P(1)(65),lamdaB => P(1)(577),lamdaOut => P(0)(65));
U_F166: entity F port map(lamdaA => P(1)(66),lamdaB => P(1)(578),lamdaOut => P(0)(66));
U_F167: entity F port map(lamdaA => P(1)(67),lamdaB => P(1)(579),lamdaOut => P(0)(67));
U_F168: entity F port map(lamdaA => P(1)(68),lamdaB => P(1)(580),lamdaOut => P(0)(68));
U_F169: entity F port map(lamdaA => P(1)(69),lamdaB => P(1)(581),lamdaOut => P(0)(69));
U_F170: entity F port map(lamdaA => P(1)(70),lamdaB => P(1)(582),lamdaOut => P(0)(70));
U_F171: entity F port map(lamdaA => P(1)(71),lamdaB => P(1)(583),lamdaOut => P(0)(71));
U_F172: entity F port map(lamdaA => P(1)(72),lamdaB => P(1)(584),lamdaOut => P(0)(72));
U_F173: entity F port map(lamdaA => P(1)(73),lamdaB => P(1)(585),lamdaOut => P(0)(73));
U_F174: entity F port map(lamdaA => P(1)(74),lamdaB => P(1)(586),lamdaOut => P(0)(74));
U_F175: entity F port map(lamdaA => P(1)(75),lamdaB => P(1)(587),lamdaOut => P(0)(75));
U_F176: entity F port map(lamdaA => P(1)(76),lamdaB => P(1)(588),lamdaOut => P(0)(76));
U_F177: entity F port map(lamdaA => P(1)(77),lamdaB => P(1)(589),lamdaOut => P(0)(77));
U_F178: entity F port map(lamdaA => P(1)(78),lamdaB => P(1)(590),lamdaOut => P(0)(78));
U_F179: entity F port map(lamdaA => P(1)(79),lamdaB => P(1)(591),lamdaOut => P(0)(79));
U_F180: entity F port map(lamdaA => P(1)(80),lamdaB => P(1)(592),lamdaOut => P(0)(80));
U_F181: entity F port map(lamdaA => P(1)(81),lamdaB => P(1)(593),lamdaOut => P(0)(81));
U_F182: entity F port map(lamdaA => P(1)(82),lamdaB => P(1)(594),lamdaOut => P(0)(82));
U_F183: entity F port map(lamdaA => P(1)(83),lamdaB => P(1)(595),lamdaOut => P(0)(83));
U_F184: entity F port map(lamdaA => P(1)(84),lamdaB => P(1)(596),lamdaOut => P(0)(84));
U_F185: entity F port map(lamdaA => P(1)(85),lamdaB => P(1)(597),lamdaOut => P(0)(85));
U_F186: entity F port map(lamdaA => P(1)(86),lamdaB => P(1)(598),lamdaOut => P(0)(86));
U_F187: entity F port map(lamdaA => P(1)(87),lamdaB => P(1)(599),lamdaOut => P(0)(87));
U_F188: entity F port map(lamdaA => P(1)(88),lamdaB => P(1)(600),lamdaOut => P(0)(88));
U_F189: entity F port map(lamdaA => P(1)(89),lamdaB => P(1)(601),lamdaOut => P(0)(89));
U_F190: entity F port map(lamdaA => P(1)(90),lamdaB => P(1)(602),lamdaOut => P(0)(90));
U_F191: entity F port map(lamdaA => P(1)(91),lamdaB => P(1)(603),lamdaOut => P(0)(91));
U_F192: entity F port map(lamdaA => P(1)(92),lamdaB => P(1)(604),lamdaOut => P(0)(92));
U_F193: entity F port map(lamdaA => P(1)(93),lamdaB => P(1)(605),lamdaOut => P(0)(93));
U_F194: entity F port map(lamdaA => P(1)(94),lamdaB => P(1)(606),lamdaOut => P(0)(94));
U_F195: entity F port map(lamdaA => P(1)(95),lamdaB => P(1)(607),lamdaOut => P(0)(95));
U_F196: entity F port map(lamdaA => P(1)(96),lamdaB => P(1)(608),lamdaOut => P(0)(96));
U_F197: entity F port map(lamdaA => P(1)(97),lamdaB => P(1)(609),lamdaOut => P(0)(97));
U_F198: entity F port map(lamdaA => P(1)(98),lamdaB => P(1)(610),lamdaOut => P(0)(98));
U_F199: entity F port map(lamdaA => P(1)(99),lamdaB => P(1)(611),lamdaOut => P(0)(99));
U_F1100: entity F port map(lamdaA => P(1)(100),lamdaB => P(1)(612),lamdaOut => P(0)(100));
U_F1101: entity F port map(lamdaA => P(1)(101),lamdaB => P(1)(613),lamdaOut => P(0)(101));
U_F1102: entity F port map(lamdaA => P(1)(102),lamdaB => P(1)(614),lamdaOut => P(0)(102));
U_F1103: entity F port map(lamdaA => P(1)(103),lamdaB => P(1)(615),lamdaOut => P(0)(103));
U_F1104: entity F port map(lamdaA => P(1)(104),lamdaB => P(1)(616),lamdaOut => P(0)(104));
U_F1105: entity F port map(lamdaA => P(1)(105),lamdaB => P(1)(617),lamdaOut => P(0)(105));
U_F1106: entity F port map(lamdaA => P(1)(106),lamdaB => P(1)(618),lamdaOut => P(0)(106));
U_F1107: entity F port map(lamdaA => P(1)(107),lamdaB => P(1)(619),lamdaOut => P(0)(107));
U_F1108: entity F port map(lamdaA => P(1)(108),lamdaB => P(1)(620),lamdaOut => P(0)(108));
U_F1109: entity F port map(lamdaA => P(1)(109),lamdaB => P(1)(621),lamdaOut => P(0)(109));
U_F1110: entity F port map(lamdaA => P(1)(110),lamdaB => P(1)(622),lamdaOut => P(0)(110));
U_F1111: entity F port map(lamdaA => P(1)(111),lamdaB => P(1)(623),lamdaOut => P(0)(111));
U_F1112: entity F port map(lamdaA => P(1)(112),lamdaB => P(1)(624),lamdaOut => P(0)(112));
U_F1113: entity F port map(lamdaA => P(1)(113),lamdaB => P(1)(625),lamdaOut => P(0)(113));
U_F1114: entity F port map(lamdaA => P(1)(114),lamdaB => P(1)(626),lamdaOut => P(0)(114));
U_F1115: entity F port map(lamdaA => P(1)(115),lamdaB => P(1)(627),lamdaOut => P(0)(115));
U_F1116: entity F port map(lamdaA => P(1)(116),lamdaB => P(1)(628),lamdaOut => P(0)(116));
U_F1117: entity F port map(lamdaA => P(1)(117),lamdaB => P(1)(629),lamdaOut => P(0)(117));
U_F1118: entity F port map(lamdaA => P(1)(118),lamdaB => P(1)(630),lamdaOut => P(0)(118));
U_F1119: entity F port map(lamdaA => P(1)(119),lamdaB => P(1)(631),lamdaOut => P(0)(119));
U_F1120: entity F port map(lamdaA => P(1)(120),lamdaB => P(1)(632),lamdaOut => P(0)(120));
U_F1121: entity F port map(lamdaA => P(1)(121),lamdaB => P(1)(633),lamdaOut => P(0)(121));
U_F1122: entity F port map(lamdaA => P(1)(122),lamdaB => P(1)(634),lamdaOut => P(0)(122));
U_F1123: entity F port map(lamdaA => P(1)(123),lamdaB => P(1)(635),lamdaOut => P(0)(123));
U_F1124: entity F port map(lamdaA => P(1)(124),lamdaB => P(1)(636),lamdaOut => P(0)(124));
U_F1125: entity F port map(lamdaA => P(1)(125),lamdaB => P(1)(637),lamdaOut => P(0)(125));
U_F1126: entity F port map(lamdaA => P(1)(126),lamdaB => P(1)(638),lamdaOut => P(0)(126));
U_F1127: entity F port map(lamdaA => P(1)(127),lamdaB => P(1)(639),lamdaOut => P(0)(127));
U_F1128: entity F port map(lamdaA => P(1)(128),lamdaB => P(1)(640),lamdaOut => P(0)(128));
U_F1129: entity F port map(lamdaA => P(1)(129),lamdaB => P(1)(641),lamdaOut => P(0)(129));
U_F1130: entity F port map(lamdaA => P(1)(130),lamdaB => P(1)(642),lamdaOut => P(0)(130));
U_F1131: entity F port map(lamdaA => P(1)(131),lamdaB => P(1)(643),lamdaOut => P(0)(131));
U_F1132: entity F port map(lamdaA => P(1)(132),lamdaB => P(1)(644),lamdaOut => P(0)(132));
U_F1133: entity F port map(lamdaA => P(1)(133),lamdaB => P(1)(645),lamdaOut => P(0)(133));
U_F1134: entity F port map(lamdaA => P(1)(134),lamdaB => P(1)(646),lamdaOut => P(0)(134));
U_F1135: entity F port map(lamdaA => P(1)(135),lamdaB => P(1)(647),lamdaOut => P(0)(135));
U_F1136: entity F port map(lamdaA => P(1)(136),lamdaB => P(1)(648),lamdaOut => P(0)(136));
U_F1137: entity F port map(lamdaA => P(1)(137),lamdaB => P(1)(649),lamdaOut => P(0)(137));
U_F1138: entity F port map(lamdaA => P(1)(138),lamdaB => P(1)(650),lamdaOut => P(0)(138));
U_F1139: entity F port map(lamdaA => P(1)(139),lamdaB => P(1)(651),lamdaOut => P(0)(139));
U_F1140: entity F port map(lamdaA => P(1)(140),lamdaB => P(1)(652),lamdaOut => P(0)(140));
U_F1141: entity F port map(lamdaA => P(1)(141),lamdaB => P(1)(653),lamdaOut => P(0)(141));
U_F1142: entity F port map(lamdaA => P(1)(142),lamdaB => P(1)(654),lamdaOut => P(0)(142));
U_F1143: entity F port map(lamdaA => P(1)(143),lamdaB => P(1)(655),lamdaOut => P(0)(143));
U_F1144: entity F port map(lamdaA => P(1)(144),lamdaB => P(1)(656),lamdaOut => P(0)(144));
U_F1145: entity F port map(lamdaA => P(1)(145),lamdaB => P(1)(657),lamdaOut => P(0)(145));
U_F1146: entity F port map(lamdaA => P(1)(146),lamdaB => P(1)(658),lamdaOut => P(0)(146));
U_F1147: entity F port map(lamdaA => P(1)(147),lamdaB => P(1)(659),lamdaOut => P(0)(147));
U_F1148: entity F port map(lamdaA => P(1)(148),lamdaB => P(1)(660),lamdaOut => P(0)(148));
U_F1149: entity F port map(lamdaA => P(1)(149),lamdaB => P(1)(661),lamdaOut => P(0)(149));
U_F1150: entity F port map(lamdaA => P(1)(150),lamdaB => P(1)(662),lamdaOut => P(0)(150));
U_F1151: entity F port map(lamdaA => P(1)(151),lamdaB => P(1)(663),lamdaOut => P(0)(151));
U_F1152: entity F port map(lamdaA => P(1)(152),lamdaB => P(1)(664),lamdaOut => P(0)(152));
U_F1153: entity F port map(lamdaA => P(1)(153),lamdaB => P(1)(665),lamdaOut => P(0)(153));
U_F1154: entity F port map(lamdaA => P(1)(154),lamdaB => P(1)(666),lamdaOut => P(0)(154));
U_F1155: entity F port map(lamdaA => P(1)(155),lamdaB => P(1)(667),lamdaOut => P(0)(155));
U_F1156: entity F port map(lamdaA => P(1)(156),lamdaB => P(1)(668),lamdaOut => P(0)(156));
U_F1157: entity F port map(lamdaA => P(1)(157),lamdaB => P(1)(669),lamdaOut => P(0)(157));
U_F1158: entity F port map(lamdaA => P(1)(158),lamdaB => P(1)(670),lamdaOut => P(0)(158));
U_F1159: entity F port map(lamdaA => P(1)(159),lamdaB => P(1)(671),lamdaOut => P(0)(159));
U_F1160: entity F port map(lamdaA => P(1)(160),lamdaB => P(1)(672),lamdaOut => P(0)(160));
U_F1161: entity F port map(lamdaA => P(1)(161),lamdaB => P(1)(673),lamdaOut => P(0)(161));
U_F1162: entity F port map(lamdaA => P(1)(162),lamdaB => P(1)(674),lamdaOut => P(0)(162));
U_F1163: entity F port map(lamdaA => P(1)(163),lamdaB => P(1)(675),lamdaOut => P(0)(163));
U_F1164: entity F port map(lamdaA => P(1)(164),lamdaB => P(1)(676),lamdaOut => P(0)(164));
U_F1165: entity F port map(lamdaA => P(1)(165),lamdaB => P(1)(677),lamdaOut => P(0)(165));
U_F1166: entity F port map(lamdaA => P(1)(166),lamdaB => P(1)(678),lamdaOut => P(0)(166));
U_F1167: entity F port map(lamdaA => P(1)(167),lamdaB => P(1)(679),lamdaOut => P(0)(167));
U_F1168: entity F port map(lamdaA => P(1)(168),lamdaB => P(1)(680),lamdaOut => P(0)(168));
U_F1169: entity F port map(lamdaA => P(1)(169),lamdaB => P(1)(681),lamdaOut => P(0)(169));
U_F1170: entity F port map(lamdaA => P(1)(170),lamdaB => P(1)(682),lamdaOut => P(0)(170));
U_F1171: entity F port map(lamdaA => P(1)(171),lamdaB => P(1)(683),lamdaOut => P(0)(171));
U_F1172: entity F port map(lamdaA => P(1)(172),lamdaB => P(1)(684),lamdaOut => P(0)(172));
U_F1173: entity F port map(lamdaA => P(1)(173),lamdaB => P(1)(685),lamdaOut => P(0)(173));
U_F1174: entity F port map(lamdaA => P(1)(174),lamdaB => P(1)(686),lamdaOut => P(0)(174));
U_F1175: entity F port map(lamdaA => P(1)(175),lamdaB => P(1)(687),lamdaOut => P(0)(175));
U_F1176: entity F port map(lamdaA => P(1)(176),lamdaB => P(1)(688),lamdaOut => P(0)(176));
U_F1177: entity F port map(lamdaA => P(1)(177),lamdaB => P(1)(689),lamdaOut => P(0)(177));
U_F1178: entity F port map(lamdaA => P(1)(178),lamdaB => P(1)(690),lamdaOut => P(0)(178));
U_F1179: entity F port map(lamdaA => P(1)(179),lamdaB => P(1)(691),lamdaOut => P(0)(179));
U_F1180: entity F port map(lamdaA => P(1)(180),lamdaB => P(1)(692),lamdaOut => P(0)(180));
U_F1181: entity F port map(lamdaA => P(1)(181),lamdaB => P(1)(693),lamdaOut => P(0)(181));
U_F1182: entity F port map(lamdaA => P(1)(182),lamdaB => P(1)(694),lamdaOut => P(0)(182));
U_F1183: entity F port map(lamdaA => P(1)(183),lamdaB => P(1)(695),lamdaOut => P(0)(183));
U_F1184: entity F port map(lamdaA => P(1)(184),lamdaB => P(1)(696),lamdaOut => P(0)(184));
U_F1185: entity F port map(lamdaA => P(1)(185),lamdaB => P(1)(697),lamdaOut => P(0)(185));
U_F1186: entity F port map(lamdaA => P(1)(186),lamdaB => P(1)(698),lamdaOut => P(0)(186));
U_F1187: entity F port map(lamdaA => P(1)(187),lamdaB => P(1)(699),lamdaOut => P(0)(187));
U_F1188: entity F port map(lamdaA => P(1)(188),lamdaB => P(1)(700),lamdaOut => P(0)(188));
U_F1189: entity F port map(lamdaA => P(1)(189),lamdaB => P(1)(701),lamdaOut => P(0)(189));
U_F1190: entity F port map(lamdaA => P(1)(190),lamdaB => P(1)(702),lamdaOut => P(0)(190));
U_F1191: entity F port map(lamdaA => P(1)(191),lamdaB => P(1)(703),lamdaOut => P(0)(191));
U_F1192: entity F port map(lamdaA => P(1)(192),lamdaB => P(1)(704),lamdaOut => P(0)(192));
U_F1193: entity F port map(lamdaA => P(1)(193),lamdaB => P(1)(705),lamdaOut => P(0)(193));
U_F1194: entity F port map(lamdaA => P(1)(194),lamdaB => P(1)(706),lamdaOut => P(0)(194));
U_F1195: entity F port map(lamdaA => P(1)(195),lamdaB => P(1)(707),lamdaOut => P(0)(195));
U_F1196: entity F port map(lamdaA => P(1)(196),lamdaB => P(1)(708),lamdaOut => P(0)(196));
U_F1197: entity F port map(lamdaA => P(1)(197),lamdaB => P(1)(709),lamdaOut => P(0)(197));
U_F1198: entity F port map(lamdaA => P(1)(198),lamdaB => P(1)(710),lamdaOut => P(0)(198));
U_F1199: entity F port map(lamdaA => P(1)(199),lamdaB => P(1)(711),lamdaOut => P(0)(199));
U_F1200: entity F port map(lamdaA => P(1)(200),lamdaB => P(1)(712),lamdaOut => P(0)(200));
U_F1201: entity F port map(lamdaA => P(1)(201),lamdaB => P(1)(713),lamdaOut => P(0)(201));
U_F1202: entity F port map(lamdaA => P(1)(202),lamdaB => P(1)(714),lamdaOut => P(0)(202));
U_F1203: entity F port map(lamdaA => P(1)(203),lamdaB => P(1)(715),lamdaOut => P(0)(203));
U_F1204: entity F port map(lamdaA => P(1)(204),lamdaB => P(1)(716),lamdaOut => P(0)(204));
U_F1205: entity F port map(lamdaA => P(1)(205),lamdaB => P(1)(717),lamdaOut => P(0)(205));
U_F1206: entity F port map(lamdaA => P(1)(206),lamdaB => P(1)(718),lamdaOut => P(0)(206));
U_F1207: entity F port map(lamdaA => P(1)(207),lamdaB => P(1)(719),lamdaOut => P(0)(207));
U_F1208: entity F port map(lamdaA => P(1)(208),lamdaB => P(1)(720),lamdaOut => P(0)(208));
U_F1209: entity F port map(lamdaA => P(1)(209),lamdaB => P(1)(721),lamdaOut => P(0)(209));
U_F1210: entity F port map(lamdaA => P(1)(210),lamdaB => P(1)(722),lamdaOut => P(0)(210));
U_F1211: entity F port map(lamdaA => P(1)(211),lamdaB => P(1)(723),lamdaOut => P(0)(211));
U_F1212: entity F port map(lamdaA => P(1)(212),lamdaB => P(1)(724),lamdaOut => P(0)(212));
U_F1213: entity F port map(lamdaA => P(1)(213),lamdaB => P(1)(725),lamdaOut => P(0)(213));
U_F1214: entity F port map(lamdaA => P(1)(214),lamdaB => P(1)(726),lamdaOut => P(0)(214));
U_F1215: entity F port map(lamdaA => P(1)(215),lamdaB => P(1)(727),lamdaOut => P(0)(215));
U_F1216: entity F port map(lamdaA => P(1)(216),lamdaB => P(1)(728),lamdaOut => P(0)(216));
U_F1217: entity F port map(lamdaA => P(1)(217),lamdaB => P(1)(729),lamdaOut => P(0)(217));
U_F1218: entity F port map(lamdaA => P(1)(218),lamdaB => P(1)(730),lamdaOut => P(0)(218));
U_F1219: entity F port map(lamdaA => P(1)(219),lamdaB => P(1)(731),lamdaOut => P(0)(219));
U_F1220: entity F port map(lamdaA => P(1)(220),lamdaB => P(1)(732),lamdaOut => P(0)(220));
U_F1221: entity F port map(lamdaA => P(1)(221),lamdaB => P(1)(733),lamdaOut => P(0)(221));
U_F1222: entity F port map(lamdaA => P(1)(222),lamdaB => P(1)(734),lamdaOut => P(0)(222));
U_F1223: entity F port map(lamdaA => P(1)(223),lamdaB => P(1)(735),lamdaOut => P(0)(223));
U_F1224: entity F port map(lamdaA => P(1)(224),lamdaB => P(1)(736),lamdaOut => P(0)(224));
U_F1225: entity F port map(lamdaA => P(1)(225),lamdaB => P(1)(737),lamdaOut => P(0)(225));
U_F1226: entity F port map(lamdaA => P(1)(226),lamdaB => P(1)(738),lamdaOut => P(0)(226));
U_F1227: entity F port map(lamdaA => P(1)(227),lamdaB => P(1)(739),lamdaOut => P(0)(227));
U_F1228: entity F port map(lamdaA => P(1)(228),lamdaB => P(1)(740),lamdaOut => P(0)(228));
U_F1229: entity F port map(lamdaA => P(1)(229),lamdaB => P(1)(741),lamdaOut => P(0)(229));
U_F1230: entity F port map(lamdaA => P(1)(230),lamdaB => P(1)(742),lamdaOut => P(0)(230));
U_F1231: entity F port map(lamdaA => P(1)(231),lamdaB => P(1)(743),lamdaOut => P(0)(231));
U_F1232: entity F port map(lamdaA => P(1)(232),lamdaB => P(1)(744),lamdaOut => P(0)(232));
U_F1233: entity F port map(lamdaA => P(1)(233),lamdaB => P(1)(745),lamdaOut => P(0)(233));
U_F1234: entity F port map(lamdaA => P(1)(234),lamdaB => P(1)(746),lamdaOut => P(0)(234));
U_F1235: entity F port map(lamdaA => P(1)(235),lamdaB => P(1)(747),lamdaOut => P(0)(235));
U_F1236: entity F port map(lamdaA => P(1)(236),lamdaB => P(1)(748),lamdaOut => P(0)(236));
U_F1237: entity F port map(lamdaA => P(1)(237),lamdaB => P(1)(749),lamdaOut => P(0)(237));
U_F1238: entity F port map(lamdaA => P(1)(238),lamdaB => P(1)(750),lamdaOut => P(0)(238));
U_F1239: entity F port map(lamdaA => P(1)(239),lamdaB => P(1)(751),lamdaOut => P(0)(239));
U_F1240: entity F port map(lamdaA => P(1)(240),lamdaB => P(1)(752),lamdaOut => P(0)(240));
U_F1241: entity F port map(lamdaA => P(1)(241),lamdaB => P(1)(753),lamdaOut => P(0)(241));
U_F1242: entity F port map(lamdaA => P(1)(242),lamdaB => P(1)(754),lamdaOut => P(0)(242));
U_F1243: entity F port map(lamdaA => P(1)(243),lamdaB => P(1)(755),lamdaOut => P(0)(243));
U_F1244: entity F port map(lamdaA => P(1)(244),lamdaB => P(1)(756),lamdaOut => P(0)(244));
U_F1245: entity F port map(lamdaA => P(1)(245),lamdaB => P(1)(757),lamdaOut => P(0)(245));
U_F1246: entity F port map(lamdaA => P(1)(246),lamdaB => P(1)(758),lamdaOut => P(0)(246));
U_F1247: entity F port map(lamdaA => P(1)(247),lamdaB => P(1)(759),lamdaOut => P(0)(247));
U_F1248: entity F port map(lamdaA => P(1)(248),lamdaB => P(1)(760),lamdaOut => P(0)(248));
U_F1249: entity F port map(lamdaA => P(1)(249),lamdaB => P(1)(761),lamdaOut => P(0)(249));
U_F1250: entity F port map(lamdaA => P(1)(250),lamdaB => P(1)(762),lamdaOut => P(0)(250));
U_F1251: entity F port map(lamdaA => P(1)(251),lamdaB => P(1)(763),lamdaOut => P(0)(251));
U_F1252: entity F port map(lamdaA => P(1)(252),lamdaB => P(1)(764),lamdaOut => P(0)(252));
U_F1253: entity F port map(lamdaA => P(1)(253),lamdaB => P(1)(765),lamdaOut => P(0)(253));
U_F1254: entity F port map(lamdaA => P(1)(254),lamdaB => P(1)(766),lamdaOut => P(0)(254));
U_F1255: entity F port map(lamdaA => P(1)(255),lamdaB => P(1)(767),lamdaOut => P(0)(255));
U_F1256: entity F port map(lamdaA => P(1)(256),lamdaB => P(1)(768),lamdaOut => P(0)(256));
U_F1257: entity F port map(lamdaA => P(1)(257),lamdaB => P(1)(769),lamdaOut => P(0)(257));
U_F1258: entity F port map(lamdaA => P(1)(258),lamdaB => P(1)(770),lamdaOut => P(0)(258));
U_F1259: entity F port map(lamdaA => P(1)(259),lamdaB => P(1)(771),lamdaOut => P(0)(259));
U_F1260: entity F port map(lamdaA => P(1)(260),lamdaB => P(1)(772),lamdaOut => P(0)(260));
U_F1261: entity F port map(lamdaA => P(1)(261),lamdaB => P(1)(773),lamdaOut => P(0)(261));
U_F1262: entity F port map(lamdaA => P(1)(262),lamdaB => P(1)(774),lamdaOut => P(0)(262));
U_F1263: entity F port map(lamdaA => P(1)(263),lamdaB => P(1)(775),lamdaOut => P(0)(263));
U_F1264: entity F port map(lamdaA => P(1)(264),lamdaB => P(1)(776),lamdaOut => P(0)(264));
U_F1265: entity F port map(lamdaA => P(1)(265),lamdaB => P(1)(777),lamdaOut => P(0)(265));
U_F1266: entity F port map(lamdaA => P(1)(266),lamdaB => P(1)(778),lamdaOut => P(0)(266));
U_F1267: entity F port map(lamdaA => P(1)(267),lamdaB => P(1)(779),lamdaOut => P(0)(267));
U_F1268: entity F port map(lamdaA => P(1)(268),lamdaB => P(1)(780),lamdaOut => P(0)(268));
U_F1269: entity F port map(lamdaA => P(1)(269),lamdaB => P(1)(781),lamdaOut => P(0)(269));
U_F1270: entity F port map(lamdaA => P(1)(270),lamdaB => P(1)(782),lamdaOut => P(0)(270));
U_F1271: entity F port map(lamdaA => P(1)(271),lamdaB => P(1)(783),lamdaOut => P(0)(271));
U_F1272: entity F port map(lamdaA => P(1)(272),lamdaB => P(1)(784),lamdaOut => P(0)(272));
U_F1273: entity F port map(lamdaA => P(1)(273),lamdaB => P(1)(785),lamdaOut => P(0)(273));
U_F1274: entity F port map(lamdaA => P(1)(274),lamdaB => P(1)(786),lamdaOut => P(0)(274));
U_F1275: entity F port map(lamdaA => P(1)(275),lamdaB => P(1)(787),lamdaOut => P(0)(275));
U_F1276: entity F port map(lamdaA => P(1)(276),lamdaB => P(1)(788),lamdaOut => P(0)(276));
U_F1277: entity F port map(lamdaA => P(1)(277),lamdaB => P(1)(789),lamdaOut => P(0)(277));
U_F1278: entity F port map(lamdaA => P(1)(278),lamdaB => P(1)(790),lamdaOut => P(0)(278));
U_F1279: entity F port map(lamdaA => P(1)(279),lamdaB => P(1)(791),lamdaOut => P(0)(279));
U_F1280: entity F port map(lamdaA => P(1)(280),lamdaB => P(1)(792),lamdaOut => P(0)(280));
U_F1281: entity F port map(lamdaA => P(1)(281),lamdaB => P(1)(793),lamdaOut => P(0)(281));
U_F1282: entity F port map(lamdaA => P(1)(282),lamdaB => P(1)(794),lamdaOut => P(0)(282));
U_F1283: entity F port map(lamdaA => P(1)(283),lamdaB => P(1)(795),lamdaOut => P(0)(283));
U_F1284: entity F port map(lamdaA => P(1)(284),lamdaB => P(1)(796),lamdaOut => P(0)(284));
U_F1285: entity F port map(lamdaA => P(1)(285),lamdaB => P(1)(797),lamdaOut => P(0)(285));
U_F1286: entity F port map(lamdaA => P(1)(286),lamdaB => P(1)(798),lamdaOut => P(0)(286));
U_F1287: entity F port map(lamdaA => P(1)(287),lamdaB => P(1)(799),lamdaOut => P(0)(287));
U_F1288: entity F port map(lamdaA => P(1)(288),lamdaB => P(1)(800),lamdaOut => P(0)(288));
U_F1289: entity F port map(lamdaA => P(1)(289),lamdaB => P(1)(801),lamdaOut => P(0)(289));
U_F1290: entity F port map(lamdaA => P(1)(290),lamdaB => P(1)(802),lamdaOut => P(0)(290));
U_F1291: entity F port map(lamdaA => P(1)(291),lamdaB => P(1)(803),lamdaOut => P(0)(291));
U_F1292: entity F port map(lamdaA => P(1)(292),lamdaB => P(1)(804),lamdaOut => P(0)(292));
U_F1293: entity F port map(lamdaA => P(1)(293),lamdaB => P(1)(805),lamdaOut => P(0)(293));
U_F1294: entity F port map(lamdaA => P(1)(294),lamdaB => P(1)(806),lamdaOut => P(0)(294));
U_F1295: entity F port map(lamdaA => P(1)(295),lamdaB => P(1)(807),lamdaOut => P(0)(295));
U_F1296: entity F port map(lamdaA => P(1)(296),lamdaB => P(1)(808),lamdaOut => P(0)(296));
U_F1297: entity F port map(lamdaA => P(1)(297),lamdaB => P(1)(809),lamdaOut => P(0)(297));
U_F1298: entity F port map(lamdaA => P(1)(298),lamdaB => P(1)(810),lamdaOut => P(0)(298));
U_F1299: entity F port map(lamdaA => P(1)(299),lamdaB => P(1)(811),lamdaOut => P(0)(299));
U_F1300: entity F port map(lamdaA => P(1)(300),lamdaB => P(1)(812),lamdaOut => P(0)(300));
U_F1301: entity F port map(lamdaA => P(1)(301),lamdaB => P(1)(813),lamdaOut => P(0)(301));
U_F1302: entity F port map(lamdaA => P(1)(302),lamdaB => P(1)(814),lamdaOut => P(0)(302));
U_F1303: entity F port map(lamdaA => P(1)(303),lamdaB => P(1)(815),lamdaOut => P(0)(303));
U_F1304: entity F port map(lamdaA => P(1)(304),lamdaB => P(1)(816),lamdaOut => P(0)(304));
U_F1305: entity F port map(lamdaA => P(1)(305),lamdaB => P(1)(817),lamdaOut => P(0)(305));
U_F1306: entity F port map(lamdaA => P(1)(306),lamdaB => P(1)(818),lamdaOut => P(0)(306));
U_F1307: entity F port map(lamdaA => P(1)(307),lamdaB => P(1)(819),lamdaOut => P(0)(307));
U_F1308: entity F port map(lamdaA => P(1)(308),lamdaB => P(1)(820),lamdaOut => P(0)(308));
U_F1309: entity F port map(lamdaA => P(1)(309),lamdaB => P(1)(821),lamdaOut => P(0)(309));
U_F1310: entity F port map(lamdaA => P(1)(310),lamdaB => P(1)(822),lamdaOut => P(0)(310));
U_F1311: entity F port map(lamdaA => P(1)(311),lamdaB => P(1)(823),lamdaOut => P(0)(311));
U_F1312: entity F port map(lamdaA => P(1)(312),lamdaB => P(1)(824),lamdaOut => P(0)(312));
U_F1313: entity F port map(lamdaA => P(1)(313),lamdaB => P(1)(825),lamdaOut => P(0)(313));
U_F1314: entity F port map(lamdaA => P(1)(314),lamdaB => P(1)(826),lamdaOut => P(0)(314));
U_F1315: entity F port map(lamdaA => P(1)(315),lamdaB => P(1)(827),lamdaOut => P(0)(315));
U_F1316: entity F port map(lamdaA => P(1)(316),lamdaB => P(1)(828),lamdaOut => P(0)(316));
U_F1317: entity F port map(lamdaA => P(1)(317),lamdaB => P(1)(829),lamdaOut => P(0)(317));
U_F1318: entity F port map(lamdaA => P(1)(318),lamdaB => P(1)(830),lamdaOut => P(0)(318));
U_F1319: entity F port map(lamdaA => P(1)(319),lamdaB => P(1)(831),lamdaOut => P(0)(319));
U_F1320: entity F port map(lamdaA => P(1)(320),lamdaB => P(1)(832),lamdaOut => P(0)(320));
U_F1321: entity F port map(lamdaA => P(1)(321),lamdaB => P(1)(833),lamdaOut => P(0)(321));
U_F1322: entity F port map(lamdaA => P(1)(322),lamdaB => P(1)(834),lamdaOut => P(0)(322));
U_F1323: entity F port map(lamdaA => P(1)(323),lamdaB => P(1)(835),lamdaOut => P(0)(323));
U_F1324: entity F port map(lamdaA => P(1)(324),lamdaB => P(1)(836),lamdaOut => P(0)(324));
U_F1325: entity F port map(lamdaA => P(1)(325),lamdaB => P(1)(837),lamdaOut => P(0)(325));
U_F1326: entity F port map(lamdaA => P(1)(326),lamdaB => P(1)(838),lamdaOut => P(0)(326));
U_F1327: entity F port map(lamdaA => P(1)(327),lamdaB => P(1)(839),lamdaOut => P(0)(327));
U_F1328: entity F port map(lamdaA => P(1)(328),lamdaB => P(1)(840),lamdaOut => P(0)(328));
U_F1329: entity F port map(lamdaA => P(1)(329),lamdaB => P(1)(841),lamdaOut => P(0)(329));
U_F1330: entity F port map(lamdaA => P(1)(330),lamdaB => P(1)(842),lamdaOut => P(0)(330));
U_F1331: entity F port map(lamdaA => P(1)(331),lamdaB => P(1)(843),lamdaOut => P(0)(331));
U_F1332: entity F port map(lamdaA => P(1)(332),lamdaB => P(1)(844),lamdaOut => P(0)(332));
U_F1333: entity F port map(lamdaA => P(1)(333),lamdaB => P(1)(845),lamdaOut => P(0)(333));
U_F1334: entity F port map(lamdaA => P(1)(334),lamdaB => P(1)(846),lamdaOut => P(0)(334));
U_F1335: entity F port map(lamdaA => P(1)(335),lamdaB => P(1)(847),lamdaOut => P(0)(335));
U_F1336: entity F port map(lamdaA => P(1)(336),lamdaB => P(1)(848),lamdaOut => P(0)(336));
U_F1337: entity F port map(lamdaA => P(1)(337),lamdaB => P(1)(849),lamdaOut => P(0)(337));
U_F1338: entity F port map(lamdaA => P(1)(338),lamdaB => P(1)(850),lamdaOut => P(0)(338));
U_F1339: entity F port map(lamdaA => P(1)(339),lamdaB => P(1)(851),lamdaOut => P(0)(339));
U_F1340: entity F port map(lamdaA => P(1)(340),lamdaB => P(1)(852),lamdaOut => P(0)(340));
U_F1341: entity F port map(lamdaA => P(1)(341),lamdaB => P(1)(853),lamdaOut => P(0)(341));
U_F1342: entity F port map(lamdaA => P(1)(342),lamdaB => P(1)(854),lamdaOut => P(0)(342));
U_F1343: entity F port map(lamdaA => P(1)(343),lamdaB => P(1)(855),lamdaOut => P(0)(343));
U_F1344: entity F port map(lamdaA => P(1)(344),lamdaB => P(1)(856),lamdaOut => P(0)(344));
U_F1345: entity F port map(lamdaA => P(1)(345),lamdaB => P(1)(857),lamdaOut => P(0)(345));
U_F1346: entity F port map(lamdaA => P(1)(346),lamdaB => P(1)(858),lamdaOut => P(0)(346));
U_F1347: entity F port map(lamdaA => P(1)(347),lamdaB => P(1)(859),lamdaOut => P(0)(347));
U_F1348: entity F port map(lamdaA => P(1)(348),lamdaB => P(1)(860),lamdaOut => P(0)(348));
U_F1349: entity F port map(lamdaA => P(1)(349),lamdaB => P(1)(861),lamdaOut => P(0)(349));
U_F1350: entity F port map(lamdaA => P(1)(350),lamdaB => P(1)(862),lamdaOut => P(0)(350));
U_F1351: entity F port map(lamdaA => P(1)(351),lamdaB => P(1)(863),lamdaOut => P(0)(351));
U_F1352: entity F port map(lamdaA => P(1)(352),lamdaB => P(1)(864),lamdaOut => P(0)(352));
U_F1353: entity F port map(lamdaA => P(1)(353),lamdaB => P(1)(865),lamdaOut => P(0)(353));
U_F1354: entity F port map(lamdaA => P(1)(354),lamdaB => P(1)(866),lamdaOut => P(0)(354));
U_F1355: entity F port map(lamdaA => P(1)(355),lamdaB => P(1)(867),lamdaOut => P(0)(355));
U_F1356: entity F port map(lamdaA => P(1)(356),lamdaB => P(1)(868),lamdaOut => P(0)(356));
U_F1357: entity F port map(lamdaA => P(1)(357),lamdaB => P(1)(869),lamdaOut => P(0)(357));
U_F1358: entity F port map(lamdaA => P(1)(358),lamdaB => P(1)(870),lamdaOut => P(0)(358));
U_F1359: entity F port map(lamdaA => P(1)(359),lamdaB => P(1)(871),lamdaOut => P(0)(359));
U_F1360: entity F port map(lamdaA => P(1)(360),lamdaB => P(1)(872),lamdaOut => P(0)(360));
U_F1361: entity F port map(lamdaA => P(1)(361),lamdaB => P(1)(873),lamdaOut => P(0)(361));
U_F1362: entity F port map(lamdaA => P(1)(362),lamdaB => P(1)(874),lamdaOut => P(0)(362));
U_F1363: entity F port map(lamdaA => P(1)(363),lamdaB => P(1)(875),lamdaOut => P(0)(363));
U_F1364: entity F port map(lamdaA => P(1)(364),lamdaB => P(1)(876),lamdaOut => P(0)(364));
U_F1365: entity F port map(lamdaA => P(1)(365),lamdaB => P(1)(877),lamdaOut => P(0)(365));
U_F1366: entity F port map(lamdaA => P(1)(366),lamdaB => P(1)(878),lamdaOut => P(0)(366));
U_F1367: entity F port map(lamdaA => P(1)(367),lamdaB => P(1)(879),lamdaOut => P(0)(367));
U_F1368: entity F port map(lamdaA => P(1)(368),lamdaB => P(1)(880),lamdaOut => P(0)(368));
U_F1369: entity F port map(lamdaA => P(1)(369),lamdaB => P(1)(881),lamdaOut => P(0)(369));
U_F1370: entity F port map(lamdaA => P(1)(370),lamdaB => P(1)(882),lamdaOut => P(0)(370));
U_F1371: entity F port map(lamdaA => P(1)(371),lamdaB => P(1)(883),lamdaOut => P(0)(371));
U_F1372: entity F port map(lamdaA => P(1)(372),lamdaB => P(1)(884),lamdaOut => P(0)(372));
U_F1373: entity F port map(lamdaA => P(1)(373),lamdaB => P(1)(885),lamdaOut => P(0)(373));
U_F1374: entity F port map(lamdaA => P(1)(374),lamdaB => P(1)(886),lamdaOut => P(0)(374));
U_F1375: entity F port map(lamdaA => P(1)(375),lamdaB => P(1)(887),lamdaOut => P(0)(375));
U_F1376: entity F port map(lamdaA => P(1)(376),lamdaB => P(1)(888),lamdaOut => P(0)(376));
U_F1377: entity F port map(lamdaA => P(1)(377),lamdaB => P(1)(889),lamdaOut => P(0)(377));
U_F1378: entity F port map(lamdaA => P(1)(378),lamdaB => P(1)(890),lamdaOut => P(0)(378));
U_F1379: entity F port map(lamdaA => P(1)(379),lamdaB => P(1)(891),lamdaOut => P(0)(379));
U_F1380: entity F port map(lamdaA => P(1)(380),lamdaB => P(1)(892),lamdaOut => P(0)(380));
U_F1381: entity F port map(lamdaA => P(1)(381),lamdaB => P(1)(893),lamdaOut => P(0)(381));
U_F1382: entity F port map(lamdaA => P(1)(382),lamdaB => P(1)(894),lamdaOut => P(0)(382));
U_F1383: entity F port map(lamdaA => P(1)(383),lamdaB => P(1)(895),lamdaOut => P(0)(383));
U_F1384: entity F port map(lamdaA => P(1)(384),lamdaB => P(1)(896),lamdaOut => P(0)(384));
U_F1385: entity F port map(lamdaA => P(1)(385),lamdaB => P(1)(897),lamdaOut => P(0)(385));
U_F1386: entity F port map(lamdaA => P(1)(386),lamdaB => P(1)(898),lamdaOut => P(0)(386));
U_F1387: entity F port map(lamdaA => P(1)(387),lamdaB => P(1)(899),lamdaOut => P(0)(387));
U_F1388: entity F port map(lamdaA => P(1)(388),lamdaB => P(1)(900),lamdaOut => P(0)(388));
U_F1389: entity F port map(lamdaA => P(1)(389),lamdaB => P(1)(901),lamdaOut => P(0)(389));
U_F1390: entity F port map(lamdaA => P(1)(390),lamdaB => P(1)(902),lamdaOut => P(0)(390));
U_F1391: entity F port map(lamdaA => P(1)(391),lamdaB => P(1)(903),lamdaOut => P(0)(391));
U_F1392: entity F port map(lamdaA => P(1)(392),lamdaB => P(1)(904),lamdaOut => P(0)(392));
U_F1393: entity F port map(lamdaA => P(1)(393),lamdaB => P(1)(905),lamdaOut => P(0)(393));
U_F1394: entity F port map(lamdaA => P(1)(394),lamdaB => P(1)(906),lamdaOut => P(0)(394));
U_F1395: entity F port map(lamdaA => P(1)(395),lamdaB => P(1)(907),lamdaOut => P(0)(395));
U_F1396: entity F port map(lamdaA => P(1)(396),lamdaB => P(1)(908),lamdaOut => P(0)(396));
U_F1397: entity F port map(lamdaA => P(1)(397),lamdaB => P(1)(909),lamdaOut => P(0)(397));
U_F1398: entity F port map(lamdaA => P(1)(398),lamdaB => P(1)(910),lamdaOut => P(0)(398));
U_F1399: entity F port map(lamdaA => P(1)(399),lamdaB => P(1)(911),lamdaOut => P(0)(399));
U_F1400: entity F port map(lamdaA => P(1)(400),lamdaB => P(1)(912),lamdaOut => P(0)(400));
U_F1401: entity F port map(lamdaA => P(1)(401),lamdaB => P(1)(913),lamdaOut => P(0)(401));
U_F1402: entity F port map(lamdaA => P(1)(402),lamdaB => P(1)(914),lamdaOut => P(0)(402));
U_F1403: entity F port map(lamdaA => P(1)(403),lamdaB => P(1)(915),lamdaOut => P(0)(403));
U_F1404: entity F port map(lamdaA => P(1)(404),lamdaB => P(1)(916),lamdaOut => P(0)(404));
U_F1405: entity F port map(lamdaA => P(1)(405),lamdaB => P(1)(917),lamdaOut => P(0)(405));
U_F1406: entity F port map(lamdaA => P(1)(406),lamdaB => P(1)(918),lamdaOut => P(0)(406));
U_F1407: entity F port map(lamdaA => P(1)(407),lamdaB => P(1)(919),lamdaOut => P(0)(407));
U_F1408: entity F port map(lamdaA => P(1)(408),lamdaB => P(1)(920),lamdaOut => P(0)(408));
U_F1409: entity F port map(lamdaA => P(1)(409),lamdaB => P(1)(921),lamdaOut => P(0)(409));
U_F1410: entity F port map(lamdaA => P(1)(410),lamdaB => P(1)(922),lamdaOut => P(0)(410));
U_F1411: entity F port map(lamdaA => P(1)(411),lamdaB => P(1)(923),lamdaOut => P(0)(411));
U_F1412: entity F port map(lamdaA => P(1)(412),lamdaB => P(1)(924),lamdaOut => P(0)(412));
U_F1413: entity F port map(lamdaA => P(1)(413),lamdaB => P(1)(925),lamdaOut => P(0)(413));
U_F1414: entity F port map(lamdaA => P(1)(414),lamdaB => P(1)(926),lamdaOut => P(0)(414));
U_F1415: entity F port map(lamdaA => P(1)(415),lamdaB => P(1)(927),lamdaOut => P(0)(415));
U_F1416: entity F port map(lamdaA => P(1)(416),lamdaB => P(1)(928),lamdaOut => P(0)(416));
U_F1417: entity F port map(lamdaA => P(1)(417),lamdaB => P(1)(929),lamdaOut => P(0)(417));
U_F1418: entity F port map(lamdaA => P(1)(418),lamdaB => P(1)(930),lamdaOut => P(0)(418));
U_F1419: entity F port map(lamdaA => P(1)(419),lamdaB => P(1)(931),lamdaOut => P(0)(419));
U_F1420: entity F port map(lamdaA => P(1)(420),lamdaB => P(1)(932),lamdaOut => P(0)(420));
U_F1421: entity F port map(lamdaA => P(1)(421),lamdaB => P(1)(933),lamdaOut => P(0)(421));
U_F1422: entity F port map(lamdaA => P(1)(422),lamdaB => P(1)(934),lamdaOut => P(0)(422));
U_F1423: entity F port map(lamdaA => P(1)(423),lamdaB => P(1)(935),lamdaOut => P(0)(423));
U_F1424: entity F port map(lamdaA => P(1)(424),lamdaB => P(1)(936),lamdaOut => P(0)(424));
U_F1425: entity F port map(lamdaA => P(1)(425),lamdaB => P(1)(937),lamdaOut => P(0)(425));
U_F1426: entity F port map(lamdaA => P(1)(426),lamdaB => P(1)(938),lamdaOut => P(0)(426));
U_F1427: entity F port map(lamdaA => P(1)(427),lamdaB => P(1)(939),lamdaOut => P(0)(427));
U_F1428: entity F port map(lamdaA => P(1)(428),lamdaB => P(1)(940),lamdaOut => P(0)(428));
U_F1429: entity F port map(lamdaA => P(1)(429),lamdaB => P(1)(941),lamdaOut => P(0)(429));
U_F1430: entity F port map(lamdaA => P(1)(430),lamdaB => P(1)(942),lamdaOut => P(0)(430));
U_F1431: entity F port map(lamdaA => P(1)(431),lamdaB => P(1)(943),lamdaOut => P(0)(431));
U_F1432: entity F port map(lamdaA => P(1)(432),lamdaB => P(1)(944),lamdaOut => P(0)(432));
U_F1433: entity F port map(lamdaA => P(1)(433),lamdaB => P(1)(945),lamdaOut => P(0)(433));
U_F1434: entity F port map(lamdaA => P(1)(434),lamdaB => P(1)(946),lamdaOut => P(0)(434));
U_F1435: entity F port map(lamdaA => P(1)(435),lamdaB => P(1)(947),lamdaOut => P(0)(435));
U_F1436: entity F port map(lamdaA => P(1)(436),lamdaB => P(1)(948),lamdaOut => P(0)(436));
U_F1437: entity F port map(lamdaA => P(1)(437),lamdaB => P(1)(949),lamdaOut => P(0)(437));
U_F1438: entity F port map(lamdaA => P(1)(438),lamdaB => P(1)(950),lamdaOut => P(0)(438));
U_F1439: entity F port map(lamdaA => P(1)(439),lamdaB => P(1)(951),lamdaOut => P(0)(439));
U_F1440: entity F port map(lamdaA => P(1)(440),lamdaB => P(1)(952),lamdaOut => P(0)(440));
U_F1441: entity F port map(lamdaA => P(1)(441),lamdaB => P(1)(953),lamdaOut => P(0)(441));
U_F1442: entity F port map(lamdaA => P(1)(442),lamdaB => P(1)(954),lamdaOut => P(0)(442));
U_F1443: entity F port map(lamdaA => P(1)(443),lamdaB => P(1)(955),lamdaOut => P(0)(443));
U_F1444: entity F port map(lamdaA => P(1)(444),lamdaB => P(1)(956),lamdaOut => P(0)(444));
U_F1445: entity F port map(lamdaA => P(1)(445),lamdaB => P(1)(957),lamdaOut => P(0)(445));
U_F1446: entity F port map(lamdaA => P(1)(446),lamdaB => P(1)(958),lamdaOut => P(0)(446));
U_F1447: entity F port map(lamdaA => P(1)(447),lamdaB => P(1)(959),lamdaOut => P(0)(447));
U_F1448: entity F port map(lamdaA => P(1)(448),lamdaB => P(1)(960),lamdaOut => P(0)(448));
U_F1449: entity F port map(lamdaA => P(1)(449),lamdaB => P(1)(961),lamdaOut => P(0)(449));
U_F1450: entity F port map(lamdaA => P(1)(450),lamdaB => P(1)(962),lamdaOut => P(0)(450));
U_F1451: entity F port map(lamdaA => P(1)(451),lamdaB => P(1)(963),lamdaOut => P(0)(451));
U_F1452: entity F port map(lamdaA => P(1)(452),lamdaB => P(1)(964),lamdaOut => P(0)(452));
U_F1453: entity F port map(lamdaA => P(1)(453),lamdaB => P(1)(965),lamdaOut => P(0)(453));
U_F1454: entity F port map(lamdaA => P(1)(454),lamdaB => P(1)(966),lamdaOut => P(0)(454));
U_F1455: entity F port map(lamdaA => P(1)(455),lamdaB => P(1)(967),lamdaOut => P(0)(455));
U_F1456: entity F port map(lamdaA => P(1)(456),lamdaB => P(1)(968),lamdaOut => P(0)(456));
U_F1457: entity F port map(lamdaA => P(1)(457),lamdaB => P(1)(969),lamdaOut => P(0)(457));
U_F1458: entity F port map(lamdaA => P(1)(458),lamdaB => P(1)(970),lamdaOut => P(0)(458));
U_F1459: entity F port map(lamdaA => P(1)(459),lamdaB => P(1)(971),lamdaOut => P(0)(459));
U_F1460: entity F port map(lamdaA => P(1)(460),lamdaB => P(1)(972),lamdaOut => P(0)(460));
U_F1461: entity F port map(lamdaA => P(1)(461),lamdaB => P(1)(973),lamdaOut => P(0)(461));
U_F1462: entity F port map(lamdaA => P(1)(462),lamdaB => P(1)(974),lamdaOut => P(0)(462));
U_F1463: entity F port map(lamdaA => P(1)(463),lamdaB => P(1)(975),lamdaOut => P(0)(463));
U_F1464: entity F port map(lamdaA => P(1)(464),lamdaB => P(1)(976),lamdaOut => P(0)(464));
U_F1465: entity F port map(lamdaA => P(1)(465),lamdaB => P(1)(977),lamdaOut => P(0)(465));
U_F1466: entity F port map(lamdaA => P(1)(466),lamdaB => P(1)(978),lamdaOut => P(0)(466));
U_F1467: entity F port map(lamdaA => P(1)(467),lamdaB => P(1)(979),lamdaOut => P(0)(467));
U_F1468: entity F port map(lamdaA => P(1)(468),lamdaB => P(1)(980),lamdaOut => P(0)(468));
U_F1469: entity F port map(lamdaA => P(1)(469),lamdaB => P(1)(981),lamdaOut => P(0)(469));
U_F1470: entity F port map(lamdaA => P(1)(470),lamdaB => P(1)(982),lamdaOut => P(0)(470));
U_F1471: entity F port map(lamdaA => P(1)(471),lamdaB => P(1)(983),lamdaOut => P(0)(471));
U_F1472: entity F port map(lamdaA => P(1)(472),lamdaB => P(1)(984),lamdaOut => P(0)(472));
U_F1473: entity F port map(lamdaA => P(1)(473),lamdaB => P(1)(985),lamdaOut => P(0)(473));
U_F1474: entity F port map(lamdaA => P(1)(474),lamdaB => P(1)(986),lamdaOut => P(0)(474));
U_F1475: entity F port map(lamdaA => P(1)(475),lamdaB => P(1)(987),lamdaOut => P(0)(475));
U_F1476: entity F port map(lamdaA => P(1)(476),lamdaB => P(1)(988),lamdaOut => P(0)(476));
U_F1477: entity F port map(lamdaA => P(1)(477),lamdaB => P(1)(989),lamdaOut => P(0)(477));
U_F1478: entity F port map(lamdaA => P(1)(478),lamdaB => P(1)(990),lamdaOut => P(0)(478));
U_F1479: entity F port map(lamdaA => P(1)(479),lamdaB => P(1)(991),lamdaOut => P(0)(479));
U_F1480: entity F port map(lamdaA => P(1)(480),lamdaB => P(1)(992),lamdaOut => P(0)(480));
U_F1481: entity F port map(lamdaA => P(1)(481),lamdaB => P(1)(993),lamdaOut => P(0)(481));
U_F1482: entity F port map(lamdaA => P(1)(482),lamdaB => P(1)(994),lamdaOut => P(0)(482));
U_F1483: entity F port map(lamdaA => P(1)(483),lamdaB => P(1)(995),lamdaOut => P(0)(483));
U_F1484: entity F port map(lamdaA => P(1)(484),lamdaB => P(1)(996),lamdaOut => P(0)(484));
U_F1485: entity F port map(lamdaA => P(1)(485),lamdaB => P(1)(997),lamdaOut => P(0)(485));
U_F1486: entity F port map(lamdaA => P(1)(486),lamdaB => P(1)(998),lamdaOut => P(0)(486));
U_F1487: entity F port map(lamdaA => P(1)(487),lamdaB => P(1)(999),lamdaOut => P(0)(487));
U_F1488: entity F port map(lamdaA => P(1)(488),lamdaB => P(1)(1000),lamdaOut => P(0)(488));
U_F1489: entity F port map(lamdaA => P(1)(489),lamdaB => P(1)(1001),lamdaOut => P(0)(489));
U_F1490: entity F port map(lamdaA => P(1)(490),lamdaB => P(1)(1002),lamdaOut => P(0)(490));
U_F1491: entity F port map(lamdaA => P(1)(491),lamdaB => P(1)(1003),lamdaOut => P(0)(491));
U_F1492: entity F port map(lamdaA => P(1)(492),lamdaB => P(1)(1004),lamdaOut => P(0)(492));
U_F1493: entity F port map(lamdaA => P(1)(493),lamdaB => P(1)(1005),lamdaOut => P(0)(493));
U_F1494: entity F port map(lamdaA => P(1)(494),lamdaB => P(1)(1006),lamdaOut => P(0)(494));
U_F1495: entity F port map(lamdaA => P(1)(495),lamdaB => P(1)(1007),lamdaOut => P(0)(495));
U_F1496: entity F port map(lamdaA => P(1)(496),lamdaB => P(1)(1008),lamdaOut => P(0)(496));
U_F1497: entity F port map(lamdaA => P(1)(497),lamdaB => P(1)(1009),lamdaOut => P(0)(497));
U_F1498: entity F port map(lamdaA => P(1)(498),lamdaB => P(1)(1010),lamdaOut => P(0)(498));
U_F1499: entity F port map(lamdaA => P(1)(499),lamdaB => P(1)(1011),lamdaOut => P(0)(499));
U_F1500: entity F port map(lamdaA => P(1)(500),lamdaB => P(1)(1012),lamdaOut => P(0)(500));
U_F1501: entity F port map(lamdaA => P(1)(501),lamdaB => P(1)(1013),lamdaOut => P(0)(501));
U_F1502: entity F port map(lamdaA => P(1)(502),lamdaB => P(1)(1014),lamdaOut => P(0)(502));
U_F1503: entity F port map(lamdaA => P(1)(503),lamdaB => P(1)(1015),lamdaOut => P(0)(503));
U_F1504: entity F port map(lamdaA => P(1)(504),lamdaB => P(1)(1016),lamdaOut => P(0)(504));
U_F1505: entity F port map(lamdaA => P(1)(505),lamdaB => P(1)(1017),lamdaOut => P(0)(505));
U_F1506: entity F port map(lamdaA => P(1)(506),lamdaB => P(1)(1018),lamdaOut => P(0)(506));
U_F1507: entity F port map(lamdaA => P(1)(507),lamdaB => P(1)(1019),lamdaOut => P(0)(507));
U_F1508: entity F port map(lamdaA => P(1)(508),lamdaB => P(1)(1020),lamdaOut => P(0)(508));
U_F1509: entity F port map(lamdaA => P(1)(509),lamdaB => P(1)(1021),lamdaOut => P(0)(509));
U_F1510: entity F port map(lamdaA => P(1)(510),lamdaB => P(1)(1022),lamdaOut => P(0)(510));
U_F1511: entity F port map(lamdaA => P(1)(511),lamdaB => P(1)(1023),lamdaOut => P(0)(511));
U_G1512: entity G port map(lamdaA => P(1)(0),lamdaB => P(1)(512),s => s(1)(0),lamdaOut => P(0)(512));
U_G1513: entity G port map(lamdaA => P(1)(1),lamdaB => P(1)(513),s => s(1)(1),lamdaOut => P(0)(513));
U_G1514: entity G port map(lamdaA => P(1)(2),lamdaB => P(1)(514),s => s(1)(2),lamdaOut => P(0)(514));
U_G1515: entity G port map(lamdaA => P(1)(3),lamdaB => P(1)(515),s => s(1)(3),lamdaOut => P(0)(515));
U_G1516: entity G port map(lamdaA => P(1)(4),lamdaB => P(1)(516),s => s(1)(4),lamdaOut => P(0)(516));
U_G1517: entity G port map(lamdaA => P(1)(5),lamdaB => P(1)(517),s => s(1)(5),lamdaOut => P(0)(517));
U_G1518: entity G port map(lamdaA => P(1)(6),lamdaB => P(1)(518),s => s(1)(6),lamdaOut => P(0)(518));
U_G1519: entity G port map(lamdaA => P(1)(7),lamdaB => P(1)(519),s => s(1)(7),lamdaOut => P(0)(519));
U_G1520: entity G port map(lamdaA => P(1)(8),lamdaB => P(1)(520),s => s(1)(8),lamdaOut => P(0)(520));
U_G1521: entity G port map(lamdaA => P(1)(9),lamdaB => P(1)(521),s => s(1)(9),lamdaOut => P(0)(521));
U_G1522: entity G port map(lamdaA => P(1)(10),lamdaB => P(1)(522),s => s(1)(10),lamdaOut => P(0)(522));
U_G1523: entity G port map(lamdaA => P(1)(11),lamdaB => P(1)(523),s => s(1)(11),lamdaOut => P(0)(523));
U_G1524: entity G port map(lamdaA => P(1)(12),lamdaB => P(1)(524),s => s(1)(12),lamdaOut => P(0)(524));
U_G1525: entity G port map(lamdaA => P(1)(13),lamdaB => P(1)(525),s => s(1)(13),lamdaOut => P(0)(525));
U_G1526: entity G port map(lamdaA => P(1)(14),lamdaB => P(1)(526),s => s(1)(14),lamdaOut => P(0)(526));
U_G1527: entity G port map(lamdaA => P(1)(15),lamdaB => P(1)(527),s => s(1)(15),lamdaOut => P(0)(527));
U_G1528: entity G port map(lamdaA => P(1)(16),lamdaB => P(1)(528),s => s(1)(16),lamdaOut => P(0)(528));
U_G1529: entity G port map(lamdaA => P(1)(17),lamdaB => P(1)(529),s => s(1)(17),lamdaOut => P(0)(529));
U_G1530: entity G port map(lamdaA => P(1)(18),lamdaB => P(1)(530),s => s(1)(18),lamdaOut => P(0)(530));
U_G1531: entity G port map(lamdaA => P(1)(19),lamdaB => P(1)(531),s => s(1)(19),lamdaOut => P(0)(531));
U_G1532: entity G port map(lamdaA => P(1)(20),lamdaB => P(1)(532),s => s(1)(20),lamdaOut => P(0)(532));
U_G1533: entity G port map(lamdaA => P(1)(21),lamdaB => P(1)(533),s => s(1)(21),lamdaOut => P(0)(533));
U_G1534: entity G port map(lamdaA => P(1)(22),lamdaB => P(1)(534),s => s(1)(22),lamdaOut => P(0)(534));
U_G1535: entity G port map(lamdaA => P(1)(23),lamdaB => P(1)(535),s => s(1)(23),lamdaOut => P(0)(535));
U_G1536: entity G port map(lamdaA => P(1)(24),lamdaB => P(1)(536),s => s(1)(24),lamdaOut => P(0)(536));
U_G1537: entity G port map(lamdaA => P(1)(25),lamdaB => P(1)(537),s => s(1)(25),lamdaOut => P(0)(537));
U_G1538: entity G port map(lamdaA => P(1)(26),lamdaB => P(1)(538),s => s(1)(26),lamdaOut => P(0)(538));
U_G1539: entity G port map(lamdaA => P(1)(27),lamdaB => P(1)(539),s => s(1)(27),lamdaOut => P(0)(539));
U_G1540: entity G port map(lamdaA => P(1)(28),lamdaB => P(1)(540),s => s(1)(28),lamdaOut => P(0)(540));
U_G1541: entity G port map(lamdaA => P(1)(29),lamdaB => P(1)(541),s => s(1)(29),lamdaOut => P(0)(541));
U_G1542: entity G port map(lamdaA => P(1)(30),lamdaB => P(1)(542),s => s(1)(30),lamdaOut => P(0)(542));
U_G1543: entity G port map(lamdaA => P(1)(31),lamdaB => P(1)(543),s => s(1)(31),lamdaOut => P(0)(543));
U_G1544: entity G port map(lamdaA => P(1)(32),lamdaB => P(1)(544),s => s(1)(32),lamdaOut => P(0)(544));
U_G1545: entity G port map(lamdaA => P(1)(33),lamdaB => P(1)(545),s => s(1)(33),lamdaOut => P(0)(545));
U_G1546: entity G port map(lamdaA => P(1)(34),lamdaB => P(1)(546),s => s(1)(34),lamdaOut => P(0)(546));
U_G1547: entity G port map(lamdaA => P(1)(35),lamdaB => P(1)(547),s => s(1)(35),lamdaOut => P(0)(547));
U_G1548: entity G port map(lamdaA => P(1)(36),lamdaB => P(1)(548),s => s(1)(36),lamdaOut => P(0)(548));
U_G1549: entity G port map(lamdaA => P(1)(37),lamdaB => P(1)(549),s => s(1)(37),lamdaOut => P(0)(549));
U_G1550: entity G port map(lamdaA => P(1)(38),lamdaB => P(1)(550),s => s(1)(38),lamdaOut => P(0)(550));
U_G1551: entity G port map(lamdaA => P(1)(39),lamdaB => P(1)(551),s => s(1)(39),lamdaOut => P(0)(551));
U_G1552: entity G port map(lamdaA => P(1)(40),lamdaB => P(1)(552),s => s(1)(40),lamdaOut => P(0)(552));
U_G1553: entity G port map(lamdaA => P(1)(41),lamdaB => P(1)(553),s => s(1)(41),lamdaOut => P(0)(553));
U_G1554: entity G port map(lamdaA => P(1)(42),lamdaB => P(1)(554),s => s(1)(42),lamdaOut => P(0)(554));
U_G1555: entity G port map(lamdaA => P(1)(43),lamdaB => P(1)(555),s => s(1)(43),lamdaOut => P(0)(555));
U_G1556: entity G port map(lamdaA => P(1)(44),lamdaB => P(1)(556),s => s(1)(44),lamdaOut => P(0)(556));
U_G1557: entity G port map(lamdaA => P(1)(45),lamdaB => P(1)(557),s => s(1)(45),lamdaOut => P(0)(557));
U_G1558: entity G port map(lamdaA => P(1)(46),lamdaB => P(1)(558),s => s(1)(46),lamdaOut => P(0)(558));
U_G1559: entity G port map(lamdaA => P(1)(47),lamdaB => P(1)(559),s => s(1)(47),lamdaOut => P(0)(559));
U_G1560: entity G port map(lamdaA => P(1)(48),lamdaB => P(1)(560),s => s(1)(48),lamdaOut => P(0)(560));
U_G1561: entity G port map(lamdaA => P(1)(49),lamdaB => P(1)(561),s => s(1)(49),lamdaOut => P(0)(561));
U_G1562: entity G port map(lamdaA => P(1)(50),lamdaB => P(1)(562),s => s(1)(50),lamdaOut => P(0)(562));
U_G1563: entity G port map(lamdaA => P(1)(51),lamdaB => P(1)(563),s => s(1)(51),lamdaOut => P(0)(563));
U_G1564: entity G port map(lamdaA => P(1)(52),lamdaB => P(1)(564),s => s(1)(52),lamdaOut => P(0)(564));
U_G1565: entity G port map(lamdaA => P(1)(53),lamdaB => P(1)(565),s => s(1)(53),lamdaOut => P(0)(565));
U_G1566: entity G port map(lamdaA => P(1)(54),lamdaB => P(1)(566),s => s(1)(54),lamdaOut => P(0)(566));
U_G1567: entity G port map(lamdaA => P(1)(55),lamdaB => P(1)(567),s => s(1)(55),lamdaOut => P(0)(567));
U_G1568: entity G port map(lamdaA => P(1)(56),lamdaB => P(1)(568),s => s(1)(56),lamdaOut => P(0)(568));
U_G1569: entity G port map(lamdaA => P(1)(57),lamdaB => P(1)(569),s => s(1)(57),lamdaOut => P(0)(569));
U_G1570: entity G port map(lamdaA => P(1)(58),lamdaB => P(1)(570),s => s(1)(58),lamdaOut => P(0)(570));
U_G1571: entity G port map(lamdaA => P(1)(59),lamdaB => P(1)(571),s => s(1)(59),lamdaOut => P(0)(571));
U_G1572: entity G port map(lamdaA => P(1)(60),lamdaB => P(1)(572),s => s(1)(60),lamdaOut => P(0)(572));
U_G1573: entity G port map(lamdaA => P(1)(61),lamdaB => P(1)(573),s => s(1)(61),lamdaOut => P(0)(573));
U_G1574: entity G port map(lamdaA => P(1)(62),lamdaB => P(1)(574),s => s(1)(62),lamdaOut => P(0)(574));
U_G1575: entity G port map(lamdaA => P(1)(63),lamdaB => P(1)(575),s => s(1)(63),lamdaOut => P(0)(575));
U_G1576: entity G port map(lamdaA => P(1)(64),lamdaB => P(1)(576),s => s(1)(64),lamdaOut => P(0)(576));
U_G1577: entity G port map(lamdaA => P(1)(65),lamdaB => P(1)(577),s => s(1)(65),lamdaOut => P(0)(577));
U_G1578: entity G port map(lamdaA => P(1)(66),lamdaB => P(1)(578),s => s(1)(66),lamdaOut => P(0)(578));
U_G1579: entity G port map(lamdaA => P(1)(67),lamdaB => P(1)(579),s => s(1)(67),lamdaOut => P(0)(579));
U_G1580: entity G port map(lamdaA => P(1)(68),lamdaB => P(1)(580),s => s(1)(68),lamdaOut => P(0)(580));
U_G1581: entity G port map(lamdaA => P(1)(69),lamdaB => P(1)(581),s => s(1)(69),lamdaOut => P(0)(581));
U_G1582: entity G port map(lamdaA => P(1)(70),lamdaB => P(1)(582),s => s(1)(70),lamdaOut => P(0)(582));
U_G1583: entity G port map(lamdaA => P(1)(71),lamdaB => P(1)(583),s => s(1)(71),lamdaOut => P(0)(583));
U_G1584: entity G port map(lamdaA => P(1)(72),lamdaB => P(1)(584),s => s(1)(72),lamdaOut => P(0)(584));
U_G1585: entity G port map(lamdaA => P(1)(73),lamdaB => P(1)(585),s => s(1)(73),lamdaOut => P(0)(585));
U_G1586: entity G port map(lamdaA => P(1)(74),lamdaB => P(1)(586),s => s(1)(74),lamdaOut => P(0)(586));
U_G1587: entity G port map(lamdaA => P(1)(75),lamdaB => P(1)(587),s => s(1)(75),lamdaOut => P(0)(587));
U_G1588: entity G port map(lamdaA => P(1)(76),lamdaB => P(1)(588),s => s(1)(76),lamdaOut => P(0)(588));
U_G1589: entity G port map(lamdaA => P(1)(77),lamdaB => P(1)(589),s => s(1)(77),lamdaOut => P(0)(589));
U_G1590: entity G port map(lamdaA => P(1)(78),lamdaB => P(1)(590),s => s(1)(78),lamdaOut => P(0)(590));
U_G1591: entity G port map(lamdaA => P(1)(79),lamdaB => P(1)(591),s => s(1)(79),lamdaOut => P(0)(591));
U_G1592: entity G port map(lamdaA => P(1)(80),lamdaB => P(1)(592),s => s(1)(80),lamdaOut => P(0)(592));
U_G1593: entity G port map(lamdaA => P(1)(81),lamdaB => P(1)(593),s => s(1)(81),lamdaOut => P(0)(593));
U_G1594: entity G port map(lamdaA => P(1)(82),lamdaB => P(1)(594),s => s(1)(82),lamdaOut => P(0)(594));
U_G1595: entity G port map(lamdaA => P(1)(83),lamdaB => P(1)(595),s => s(1)(83),lamdaOut => P(0)(595));
U_G1596: entity G port map(lamdaA => P(1)(84),lamdaB => P(1)(596),s => s(1)(84),lamdaOut => P(0)(596));
U_G1597: entity G port map(lamdaA => P(1)(85),lamdaB => P(1)(597),s => s(1)(85),lamdaOut => P(0)(597));
U_G1598: entity G port map(lamdaA => P(1)(86),lamdaB => P(1)(598),s => s(1)(86),lamdaOut => P(0)(598));
U_G1599: entity G port map(lamdaA => P(1)(87),lamdaB => P(1)(599),s => s(1)(87),lamdaOut => P(0)(599));
U_G1600: entity G port map(lamdaA => P(1)(88),lamdaB => P(1)(600),s => s(1)(88),lamdaOut => P(0)(600));
U_G1601: entity G port map(lamdaA => P(1)(89),lamdaB => P(1)(601),s => s(1)(89),lamdaOut => P(0)(601));
U_G1602: entity G port map(lamdaA => P(1)(90),lamdaB => P(1)(602),s => s(1)(90),lamdaOut => P(0)(602));
U_G1603: entity G port map(lamdaA => P(1)(91),lamdaB => P(1)(603),s => s(1)(91),lamdaOut => P(0)(603));
U_G1604: entity G port map(lamdaA => P(1)(92),lamdaB => P(1)(604),s => s(1)(92),lamdaOut => P(0)(604));
U_G1605: entity G port map(lamdaA => P(1)(93),lamdaB => P(1)(605),s => s(1)(93),lamdaOut => P(0)(605));
U_G1606: entity G port map(lamdaA => P(1)(94),lamdaB => P(1)(606),s => s(1)(94),lamdaOut => P(0)(606));
U_G1607: entity G port map(lamdaA => P(1)(95),lamdaB => P(1)(607),s => s(1)(95),lamdaOut => P(0)(607));
U_G1608: entity G port map(lamdaA => P(1)(96),lamdaB => P(1)(608),s => s(1)(96),lamdaOut => P(0)(608));
U_G1609: entity G port map(lamdaA => P(1)(97),lamdaB => P(1)(609),s => s(1)(97),lamdaOut => P(0)(609));
U_G1610: entity G port map(lamdaA => P(1)(98),lamdaB => P(1)(610),s => s(1)(98),lamdaOut => P(0)(610));
U_G1611: entity G port map(lamdaA => P(1)(99),lamdaB => P(1)(611),s => s(1)(99),lamdaOut => P(0)(611));
U_G1612: entity G port map(lamdaA => P(1)(100),lamdaB => P(1)(612),s => s(1)(100),lamdaOut => P(0)(612));
U_G1613: entity G port map(lamdaA => P(1)(101),lamdaB => P(1)(613),s => s(1)(101),lamdaOut => P(0)(613));
U_G1614: entity G port map(lamdaA => P(1)(102),lamdaB => P(1)(614),s => s(1)(102),lamdaOut => P(0)(614));
U_G1615: entity G port map(lamdaA => P(1)(103),lamdaB => P(1)(615),s => s(1)(103),lamdaOut => P(0)(615));
U_G1616: entity G port map(lamdaA => P(1)(104),lamdaB => P(1)(616),s => s(1)(104),lamdaOut => P(0)(616));
U_G1617: entity G port map(lamdaA => P(1)(105),lamdaB => P(1)(617),s => s(1)(105),lamdaOut => P(0)(617));
U_G1618: entity G port map(lamdaA => P(1)(106),lamdaB => P(1)(618),s => s(1)(106),lamdaOut => P(0)(618));
U_G1619: entity G port map(lamdaA => P(1)(107),lamdaB => P(1)(619),s => s(1)(107),lamdaOut => P(0)(619));
U_G1620: entity G port map(lamdaA => P(1)(108),lamdaB => P(1)(620),s => s(1)(108),lamdaOut => P(0)(620));
U_G1621: entity G port map(lamdaA => P(1)(109),lamdaB => P(1)(621),s => s(1)(109),lamdaOut => P(0)(621));
U_G1622: entity G port map(lamdaA => P(1)(110),lamdaB => P(1)(622),s => s(1)(110),lamdaOut => P(0)(622));
U_G1623: entity G port map(lamdaA => P(1)(111),lamdaB => P(1)(623),s => s(1)(111),lamdaOut => P(0)(623));
U_G1624: entity G port map(lamdaA => P(1)(112),lamdaB => P(1)(624),s => s(1)(112),lamdaOut => P(0)(624));
U_G1625: entity G port map(lamdaA => P(1)(113),lamdaB => P(1)(625),s => s(1)(113),lamdaOut => P(0)(625));
U_G1626: entity G port map(lamdaA => P(1)(114),lamdaB => P(1)(626),s => s(1)(114),lamdaOut => P(0)(626));
U_G1627: entity G port map(lamdaA => P(1)(115),lamdaB => P(1)(627),s => s(1)(115),lamdaOut => P(0)(627));
U_G1628: entity G port map(lamdaA => P(1)(116),lamdaB => P(1)(628),s => s(1)(116),lamdaOut => P(0)(628));
U_G1629: entity G port map(lamdaA => P(1)(117),lamdaB => P(1)(629),s => s(1)(117),lamdaOut => P(0)(629));
U_G1630: entity G port map(lamdaA => P(1)(118),lamdaB => P(1)(630),s => s(1)(118),lamdaOut => P(0)(630));
U_G1631: entity G port map(lamdaA => P(1)(119),lamdaB => P(1)(631),s => s(1)(119),lamdaOut => P(0)(631));
U_G1632: entity G port map(lamdaA => P(1)(120),lamdaB => P(1)(632),s => s(1)(120),lamdaOut => P(0)(632));
U_G1633: entity G port map(lamdaA => P(1)(121),lamdaB => P(1)(633),s => s(1)(121),lamdaOut => P(0)(633));
U_G1634: entity G port map(lamdaA => P(1)(122),lamdaB => P(1)(634),s => s(1)(122),lamdaOut => P(0)(634));
U_G1635: entity G port map(lamdaA => P(1)(123),lamdaB => P(1)(635),s => s(1)(123),lamdaOut => P(0)(635));
U_G1636: entity G port map(lamdaA => P(1)(124),lamdaB => P(1)(636),s => s(1)(124),lamdaOut => P(0)(636));
U_G1637: entity G port map(lamdaA => P(1)(125),lamdaB => P(1)(637),s => s(1)(125),lamdaOut => P(0)(637));
U_G1638: entity G port map(lamdaA => P(1)(126),lamdaB => P(1)(638),s => s(1)(126),lamdaOut => P(0)(638));
U_G1639: entity G port map(lamdaA => P(1)(127),lamdaB => P(1)(639),s => s(1)(127),lamdaOut => P(0)(639));
U_G1640: entity G port map(lamdaA => P(1)(128),lamdaB => P(1)(640),s => s(1)(128),lamdaOut => P(0)(640));
U_G1641: entity G port map(lamdaA => P(1)(129),lamdaB => P(1)(641),s => s(1)(129),lamdaOut => P(0)(641));
U_G1642: entity G port map(lamdaA => P(1)(130),lamdaB => P(1)(642),s => s(1)(130),lamdaOut => P(0)(642));
U_G1643: entity G port map(lamdaA => P(1)(131),lamdaB => P(1)(643),s => s(1)(131),lamdaOut => P(0)(643));
U_G1644: entity G port map(lamdaA => P(1)(132),lamdaB => P(1)(644),s => s(1)(132),lamdaOut => P(0)(644));
U_G1645: entity G port map(lamdaA => P(1)(133),lamdaB => P(1)(645),s => s(1)(133),lamdaOut => P(0)(645));
U_G1646: entity G port map(lamdaA => P(1)(134),lamdaB => P(1)(646),s => s(1)(134),lamdaOut => P(0)(646));
U_G1647: entity G port map(lamdaA => P(1)(135),lamdaB => P(1)(647),s => s(1)(135),lamdaOut => P(0)(647));
U_G1648: entity G port map(lamdaA => P(1)(136),lamdaB => P(1)(648),s => s(1)(136),lamdaOut => P(0)(648));
U_G1649: entity G port map(lamdaA => P(1)(137),lamdaB => P(1)(649),s => s(1)(137),lamdaOut => P(0)(649));
U_G1650: entity G port map(lamdaA => P(1)(138),lamdaB => P(1)(650),s => s(1)(138),lamdaOut => P(0)(650));
U_G1651: entity G port map(lamdaA => P(1)(139),lamdaB => P(1)(651),s => s(1)(139),lamdaOut => P(0)(651));
U_G1652: entity G port map(lamdaA => P(1)(140),lamdaB => P(1)(652),s => s(1)(140),lamdaOut => P(0)(652));
U_G1653: entity G port map(lamdaA => P(1)(141),lamdaB => P(1)(653),s => s(1)(141),lamdaOut => P(0)(653));
U_G1654: entity G port map(lamdaA => P(1)(142),lamdaB => P(1)(654),s => s(1)(142),lamdaOut => P(0)(654));
U_G1655: entity G port map(lamdaA => P(1)(143),lamdaB => P(1)(655),s => s(1)(143),lamdaOut => P(0)(655));
U_G1656: entity G port map(lamdaA => P(1)(144),lamdaB => P(1)(656),s => s(1)(144),lamdaOut => P(0)(656));
U_G1657: entity G port map(lamdaA => P(1)(145),lamdaB => P(1)(657),s => s(1)(145),lamdaOut => P(0)(657));
U_G1658: entity G port map(lamdaA => P(1)(146),lamdaB => P(1)(658),s => s(1)(146),lamdaOut => P(0)(658));
U_G1659: entity G port map(lamdaA => P(1)(147),lamdaB => P(1)(659),s => s(1)(147),lamdaOut => P(0)(659));
U_G1660: entity G port map(lamdaA => P(1)(148),lamdaB => P(1)(660),s => s(1)(148),lamdaOut => P(0)(660));
U_G1661: entity G port map(lamdaA => P(1)(149),lamdaB => P(1)(661),s => s(1)(149),lamdaOut => P(0)(661));
U_G1662: entity G port map(lamdaA => P(1)(150),lamdaB => P(1)(662),s => s(1)(150),lamdaOut => P(0)(662));
U_G1663: entity G port map(lamdaA => P(1)(151),lamdaB => P(1)(663),s => s(1)(151),lamdaOut => P(0)(663));
U_G1664: entity G port map(lamdaA => P(1)(152),lamdaB => P(1)(664),s => s(1)(152),lamdaOut => P(0)(664));
U_G1665: entity G port map(lamdaA => P(1)(153),lamdaB => P(1)(665),s => s(1)(153),lamdaOut => P(0)(665));
U_G1666: entity G port map(lamdaA => P(1)(154),lamdaB => P(1)(666),s => s(1)(154),lamdaOut => P(0)(666));
U_G1667: entity G port map(lamdaA => P(1)(155),lamdaB => P(1)(667),s => s(1)(155),lamdaOut => P(0)(667));
U_G1668: entity G port map(lamdaA => P(1)(156),lamdaB => P(1)(668),s => s(1)(156),lamdaOut => P(0)(668));
U_G1669: entity G port map(lamdaA => P(1)(157),lamdaB => P(1)(669),s => s(1)(157),lamdaOut => P(0)(669));
U_G1670: entity G port map(lamdaA => P(1)(158),lamdaB => P(1)(670),s => s(1)(158),lamdaOut => P(0)(670));
U_G1671: entity G port map(lamdaA => P(1)(159),lamdaB => P(1)(671),s => s(1)(159),lamdaOut => P(0)(671));
U_G1672: entity G port map(lamdaA => P(1)(160),lamdaB => P(1)(672),s => s(1)(160),lamdaOut => P(0)(672));
U_G1673: entity G port map(lamdaA => P(1)(161),lamdaB => P(1)(673),s => s(1)(161),lamdaOut => P(0)(673));
U_G1674: entity G port map(lamdaA => P(1)(162),lamdaB => P(1)(674),s => s(1)(162),lamdaOut => P(0)(674));
U_G1675: entity G port map(lamdaA => P(1)(163),lamdaB => P(1)(675),s => s(1)(163),lamdaOut => P(0)(675));
U_G1676: entity G port map(lamdaA => P(1)(164),lamdaB => P(1)(676),s => s(1)(164),lamdaOut => P(0)(676));
U_G1677: entity G port map(lamdaA => P(1)(165),lamdaB => P(1)(677),s => s(1)(165),lamdaOut => P(0)(677));
U_G1678: entity G port map(lamdaA => P(1)(166),lamdaB => P(1)(678),s => s(1)(166),lamdaOut => P(0)(678));
U_G1679: entity G port map(lamdaA => P(1)(167),lamdaB => P(1)(679),s => s(1)(167),lamdaOut => P(0)(679));
U_G1680: entity G port map(lamdaA => P(1)(168),lamdaB => P(1)(680),s => s(1)(168),lamdaOut => P(0)(680));
U_G1681: entity G port map(lamdaA => P(1)(169),lamdaB => P(1)(681),s => s(1)(169),lamdaOut => P(0)(681));
U_G1682: entity G port map(lamdaA => P(1)(170),lamdaB => P(1)(682),s => s(1)(170),lamdaOut => P(0)(682));
U_G1683: entity G port map(lamdaA => P(1)(171),lamdaB => P(1)(683),s => s(1)(171),lamdaOut => P(0)(683));
U_G1684: entity G port map(lamdaA => P(1)(172),lamdaB => P(1)(684),s => s(1)(172),lamdaOut => P(0)(684));
U_G1685: entity G port map(lamdaA => P(1)(173),lamdaB => P(1)(685),s => s(1)(173),lamdaOut => P(0)(685));
U_G1686: entity G port map(lamdaA => P(1)(174),lamdaB => P(1)(686),s => s(1)(174),lamdaOut => P(0)(686));
U_G1687: entity G port map(lamdaA => P(1)(175),lamdaB => P(1)(687),s => s(1)(175),lamdaOut => P(0)(687));
U_G1688: entity G port map(lamdaA => P(1)(176),lamdaB => P(1)(688),s => s(1)(176),lamdaOut => P(0)(688));
U_G1689: entity G port map(lamdaA => P(1)(177),lamdaB => P(1)(689),s => s(1)(177),lamdaOut => P(0)(689));
U_G1690: entity G port map(lamdaA => P(1)(178),lamdaB => P(1)(690),s => s(1)(178),lamdaOut => P(0)(690));
U_G1691: entity G port map(lamdaA => P(1)(179),lamdaB => P(1)(691),s => s(1)(179),lamdaOut => P(0)(691));
U_G1692: entity G port map(lamdaA => P(1)(180),lamdaB => P(1)(692),s => s(1)(180),lamdaOut => P(0)(692));
U_G1693: entity G port map(lamdaA => P(1)(181),lamdaB => P(1)(693),s => s(1)(181),lamdaOut => P(0)(693));
U_G1694: entity G port map(lamdaA => P(1)(182),lamdaB => P(1)(694),s => s(1)(182),lamdaOut => P(0)(694));
U_G1695: entity G port map(lamdaA => P(1)(183),lamdaB => P(1)(695),s => s(1)(183),lamdaOut => P(0)(695));
U_G1696: entity G port map(lamdaA => P(1)(184),lamdaB => P(1)(696),s => s(1)(184),lamdaOut => P(0)(696));
U_G1697: entity G port map(lamdaA => P(1)(185),lamdaB => P(1)(697),s => s(1)(185),lamdaOut => P(0)(697));
U_G1698: entity G port map(lamdaA => P(1)(186),lamdaB => P(1)(698),s => s(1)(186),lamdaOut => P(0)(698));
U_G1699: entity G port map(lamdaA => P(1)(187),lamdaB => P(1)(699),s => s(1)(187),lamdaOut => P(0)(699));
U_G1700: entity G port map(lamdaA => P(1)(188),lamdaB => P(1)(700),s => s(1)(188),lamdaOut => P(0)(700));
U_G1701: entity G port map(lamdaA => P(1)(189),lamdaB => P(1)(701),s => s(1)(189),lamdaOut => P(0)(701));
U_G1702: entity G port map(lamdaA => P(1)(190),lamdaB => P(1)(702),s => s(1)(190),lamdaOut => P(0)(702));
U_G1703: entity G port map(lamdaA => P(1)(191),lamdaB => P(1)(703),s => s(1)(191),lamdaOut => P(0)(703));
U_G1704: entity G port map(lamdaA => P(1)(192),lamdaB => P(1)(704),s => s(1)(192),lamdaOut => P(0)(704));
U_G1705: entity G port map(lamdaA => P(1)(193),lamdaB => P(1)(705),s => s(1)(193),lamdaOut => P(0)(705));
U_G1706: entity G port map(lamdaA => P(1)(194),lamdaB => P(1)(706),s => s(1)(194),lamdaOut => P(0)(706));
U_G1707: entity G port map(lamdaA => P(1)(195),lamdaB => P(1)(707),s => s(1)(195),lamdaOut => P(0)(707));
U_G1708: entity G port map(lamdaA => P(1)(196),lamdaB => P(1)(708),s => s(1)(196),lamdaOut => P(0)(708));
U_G1709: entity G port map(lamdaA => P(1)(197),lamdaB => P(1)(709),s => s(1)(197),lamdaOut => P(0)(709));
U_G1710: entity G port map(lamdaA => P(1)(198),lamdaB => P(1)(710),s => s(1)(198),lamdaOut => P(0)(710));
U_G1711: entity G port map(lamdaA => P(1)(199),lamdaB => P(1)(711),s => s(1)(199),lamdaOut => P(0)(711));
U_G1712: entity G port map(lamdaA => P(1)(200),lamdaB => P(1)(712),s => s(1)(200),lamdaOut => P(0)(712));
U_G1713: entity G port map(lamdaA => P(1)(201),lamdaB => P(1)(713),s => s(1)(201),lamdaOut => P(0)(713));
U_G1714: entity G port map(lamdaA => P(1)(202),lamdaB => P(1)(714),s => s(1)(202),lamdaOut => P(0)(714));
U_G1715: entity G port map(lamdaA => P(1)(203),lamdaB => P(1)(715),s => s(1)(203),lamdaOut => P(0)(715));
U_G1716: entity G port map(lamdaA => P(1)(204),lamdaB => P(1)(716),s => s(1)(204),lamdaOut => P(0)(716));
U_G1717: entity G port map(lamdaA => P(1)(205),lamdaB => P(1)(717),s => s(1)(205),lamdaOut => P(0)(717));
U_G1718: entity G port map(lamdaA => P(1)(206),lamdaB => P(1)(718),s => s(1)(206),lamdaOut => P(0)(718));
U_G1719: entity G port map(lamdaA => P(1)(207),lamdaB => P(1)(719),s => s(1)(207),lamdaOut => P(0)(719));
U_G1720: entity G port map(lamdaA => P(1)(208),lamdaB => P(1)(720),s => s(1)(208),lamdaOut => P(0)(720));
U_G1721: entity G port map(lamdaA => P(1)(209),lamdaB => P(1)(721),s => s(1)(209),lamdaOut => P(0)(721));
U_G1722: entity G port map(lamdaA => P(1)(210),lamdaB => P(1)(722),s => s(1)(210),lamdaOut => P(0)(722));
U_G1723: entity G port map(lamdaA => P(1)(211),lamdaB => P(1)(723),s => s(1)(211),lamdaOut => P(0)(723));
U_G1724: entity G port map(lamdaA => P(1)(212),lamdaB => P(1)(724),s => s(1)(212),lamdaOut => P(0)(724));
U_G1725: entity G port map(lamdaA => P(1)(213),lamdaB => P(1)(725),s => s(1)(213),lamdaOut => P(0)(725));
U_G1726: entity G port map(lamdaA => P(1)(214),lamdaB => P(1)(726),s => s(1)(214),lamdaOut => P(0)(726));
U_G1727: entity G port map(lamdaA => P(1)(215),lamdaB => P(1)(727),s => s(1)(215),lamdaOut => P(0)(727));
U_G1728: entity G port map(lamdaA => P(1)(216),lamdaB => P(1)(728),s => s(1)(216),lamdaOut => P(0)(728));
U_G1729: entity G port map(lamdaA => P(1)(217),lamdaB => P(1)(729),s => s(1)(217),lamdaOut => P(0)(729));
U_G1730: entity G port map(lamdaA => P(1)(218),lamdaB => P(1)(730),s => s(1)(218),lamdaOut => P(0)(730));
U_G1731: entity G port map(lamdaA => P(1)(219),lamdaB => P(1)(731),s => s(1)(219),lamdaOut => P(0)(731));
U_G1732: entity G port map(lamdaA => P(1)(220),lamdaB => P(1)(732),s => s(1)(220),lamdaOut => P(0)(732));
U_G1733: entity G port map(lamdaA => P(1)(221),lamdaB => P(1)(733),s => s(1)(221),lamdaOut => P(0)(733));
U_G1734: entity G port map(lamdaA => P(1)(222),lamdaB => P(1)(734),s => s(1)(222),lamdaOut => P(0)(734));
U_G1735: entity G port map(lamdaA => P(1)(223),lamdaB => P(1)(735),s => s(1)(223),lamdaOut => P(0)(735));
U_G1736: entity G port map(lamdaA => P(1)(224),lamdaB => P(1)(736),s => s(1)(224),lamdaOut => P(0)(736));
U_G1737: entity G port map(lamdaA => P(1)(225),lamdaB => P(1)(737),s => s(1)(225),lamdaOut => P(0)(737));
U_G1738: entity G port map(lamdaA => P(1)(226),lamdaB => P(1)(738),s => s(1)(226),lamdaOut => P(0)(738));
U_G1739: entity G port map(lamdaA => P(1)(227),lamdaB => P(1)(739),s => s(1)(227),lamdaOut => P(0)(739));
U_G1740: entity G port map(lamdaA => P(1)(228),lamdaB => P(1)(740),s => s(1)(228),lamdaOut => P(0)(740));
U_G1741: entity G port map(lamdaA => P(1)(229),lamdaB => P(1)(741),s => s(1)(229),lamdaOut => P(0)(741));
U_G1742: entity G port map(lamdaA => P(1)(230),lamdaB => P(1)(742),s => s(1)(230),lamdaOut => P(0)(742));
U_G1743: entity G port map(lamdaA => P(1)(231),lamdaB => P(1)(743),s => s(1)(231),lamdaOut => P(0)(743));
U_G1744: entity G port map(lamdaA => P(1)(232),lamdaB => P(1)(744),s => s(1)(232),lamdaOut => P(0)(744));
U_G1745: entity G port map(lamdaA => P(1)(233),lamdaB => P(1)(745),s => s(1)(233),lamdaOut => P(0)(745));
U_G1746: entity G port map(lamdaA => P(1)(234),lamdaB => P(1)(746),s => s(1)(234),lamdaOut => P(0)(746));
U_G1747: entity G port map(lamdaA => P(1)(235),lamdaB => P(1)(747),s => s(1)(235),lamdaOut => P(0)(747));
U_G1748: entity G port map(lamdaA => P(1)(236),lamdaB => P(1)(748),s => s(1)(236),lamdaOut => P(0)(748));
U_G1749: entity G port map(lamdaA => P(1)(237),lamdaB => P(1)(749),s => s(1)(237),lamdaOut => P(0)(749));
U_G1750: entity G port map(lamdaA => P(1)(238),lamdaB => P(1)(750),s => s(1)(238),lamdaOut => P(0)(750));
U_G1751: entity G port map(lamdaA => P(1)(239),lamdaB => P(1)(751),s => s(1)(239),lamdaOut => P(0)(751));
U_G1752: entity G port map(lamdaA => P(1)(240),lamdaB => P(1)(752),s => s(1)(240),lamdaOut => P(0)(752));
U_G1753: entity G port map(lamdaA => P(1)(241),lamdaB => P(1)(753),s => s(1)(241),lamdaOut => P(0)(753));
U_G1754: entity G port map(lamdaA => P(1)(242),lamdaB => P(1)(754),s => s(1)(242),lamdaOut => P(0)(754));
U_G1755: entity G port map(lamdaA => P(1)(243),lamdaB => P(1)(755),s => s(1)(243),lamdaOut => P(0)(755));
U_G1756: entity G port map(lamdaA => P(1)(244),lamdaB => P(1)(756),s => s(1)(244),lamdaOut => P(0)(756));
U_G1757: entity G port map(lamdaA => P(1)(245),lamdaB => P(1)(757),s => s(1)(245),lamdaOut => P(0)(757));
U_G1758: entity G port map(lamdaA => P(1)(246),lamdaB => P(1)(758),s => s(1)(246),lamdaOut => P(0)(758));
U_G1759: entity G port map(lamdaA => P(1)(247),lamdaB => P(1)(759),s => s(1)(247),lamdaOut => P(0)(759));
U_G1760: entity G port map(lamdaA => P(1)(248),lamdaB => P(1)(760),s => s(1)(248),lamdaOut => P(0)(760));
U_G1761: entity G port map(lamdaA => P(1)(249),lamdaB => P(1)(761),s => s(1)(249),lamdaOut => P(0)(761));
U_G1762: entity G port map(lamdaA => P(1)(250),lamdaB => P(1)(762),s => s(1)(250),lamdaOut => P(0)(762));
U_G1763: entity G port map(lamdaA => P(1)(251),lamdaB => P(1)(763),s => s(1)(251),lamdaOut => P(0)(763));
U_G1764: entity G port map(lamdaA => P(1)(252),lamdaB => P(1)(764),s => s(1)(252),lamdaOut => P(0)(764));
U_G1765: entity G port map(lamdaA => P(1)(253),lamdaB => P(1)(765),s => s(1)(253),lamdaOut => P(0)(765));
U_G1766: entity G port map(lamdaA => P(1)(254),lamdaB => P(1)(766),s => s(1)(254),lamdaOut => P(0)(766));
U_G1767: entity G port map(lamdaA => P(1)(255),lamdaB => P(1)(767),s => s(1)(255),lamdaOut => P(0)(767));
U_G1768: entity G port map(lamdaA => P(1)(256),lamdaB => P(1)(768),s => s(1)(256),lamdaOut => P(0)(768));
U_G1769: entity G port map(lamdaA => P(1)(257),lamdaB => P(1)(769),s => s(1)(257),lamdaOut => P(0)(769));
U_G1770: entity G port map(lamdaA => P(1)(258),lamdaB => P(1)(770),s => s(1)(258),lamdaOut => P(0)(770));
U_G1771: entity G port map(lamdaA => P(1)(259),lamdaB => P(1)(771),s => s(1)(259),lamdaOut => P(0)(771));
U_G1772: entity G port map(lamdaA => P(1)(260),lamdaB => P(1)(772),s => s(1)(260),lamdaOut => P(0)(772));
U_G1773: entity G port map(lamdaA => P(1)(261),lamdaB => P(1)(773),s => s(1)(261),lamdaOut => P(0)(773));
U_G1774: entity G port map(lamdaA => P(1)(262),lamdaB => P(1)(774),s => s(1)(262),lamdaOut => P(0)(774));
U_G1775: entity G port map(lamdaA => P(1)(263),lamdaB => P(1)(775),s => s(1)(263),lamdaOut => P(0)(775));
U_G1776: entity G port map(lamdaA => P(1)(264),lamdaB => P(1)(776),s => s(1)(264),lamdaOut => P(0)(776));
U_G1777: entity G port map(lamdaA => P(1)(265),lamdaB => P(1)(777),s => s(1)(265),lamdaOut => P(0)(777));
U_G1778: entity G port map(lamdaA => P(1)(266),lamdaB => P(1)(778),s => s(1)(266),lamdaOut => P(0)(778));
U_G1779: entity G port map(lamdaA => P(1)(267),lamdaB => P(1)(779),s => s(1)(267),lamdaOut => P(0)(779));
U_G1780: entity G port map(lamdaA => P(1)(268),lamdaB => P(1)(780),s => s(1)(268),lamdaOut => P(0)(780));
U_G1781: entity G port map(lamdaA => P(1)(269),lamdaB => P(1)(781),s => s(1)(269),lamdaOut => P(0)(781));
U_G1782: entity G port map(lamdaA => P(1)(270),lamdaB => P(1)(782),s => s(1)(270),lamdaOut => P(0)(782));
U_G1783: entity G port map(lamdaA => P(1)(271),lamdaB => P(1)(783),s => s(1)(271),lamdaOut => P(0)(783));
U_G1784: entity G port map(lamdaA => P(1)(272),lamdaB => P(1)(784),s => s(1)(272),lamdaOut => P(0)(784));
U_G1785: entity G port map(lamdaA => P(1)(273),lamdaB => P(1)(785),s => s(1)(273),lamdaOut => P(0)(785));
U_G1786: entity G port map(lamdaA => P(1)(274),lamdaB => P(1)(786),s => s(1)(274),lamdaOut => P(0)(786));
U_G1787: entity G port map(lamdaA => P(1)(275),lamdaB => P(1)(787),s => s(1)(275),lamdaOut => P(0)(787));
U_G1788: entity G port map(lamdaA => P(1)(276),lamdaB => P(1)(788),s => s(1)(276),lamdaOut => P(0)(788));
U_G1789: entity G port map(lamdaA => P(1)(277),lamdaB => P(1)(789),s => s(1)(277),lamdaOut => P(0)(789));
U_G1790: entity G port map(lamdaA => P(1)(278),lamdaB => P(1)(790),s => s(1)(278),lamdaOut => P(0)(790));
U_G1791: entity G port map(lamdaA => P(1)(279),lamdaB => P(1)(791),s => s(1)(279),lamdaOut => P(0)(791));
U_G1792: entity G port map(lamdaA => P(1)(280),lamdaB => P(1)(792),s => s(1)(280),lamdaOut => P(0)(792));
U_G1793: entity G port map(lamdaA => P(1)(281),lamdaB => P(1)(793),s => s(1)(281),lamdaOut => P(0)(793));
U_G1794: entity G port map(lamdaA => P(1)(282),lamdaB => P(1)(794),s => s(1)(282),lamdaOut => P(0)(794));
U_G1795: entity G port map(lamdaA => P(1)(283),lamdaB => P(1)(795),s => s(1)(283),lamdaOut => P(0)(795));
U_G1796: entity G port map(lamdaA => P(1)(284),lamdaB => P(1)(796),s => s(1)(284),lamdaOut => P(0)(796));
U_G1797: entity G port map(lamdaA => P(1)(285),lamdaB => P(1)(797),s => s(1)(285),lamdaOut => P(0)(797));
U_G1798: entity G port map(lamdaA => P(1)(286),lamdaB => P(1)(798),s => s(1)(286),lamdaOut => P(0)(798));
U_G1799: entity G port map(lamdaA => P(1)(287),lamdaB => P(1)(799),s => s(1)(287),lamdaOut => P(0)(799));
U_G1800: entity G port map(lamdaA => P(1)(288),lamdaB => P(1)(800),s => s(1)(288),lamdaOut => P(0)(800));
U_G1801: entity G port map(lamdaA => P(1)(289),lamdaB => P(1)(801),s => s(1)(289),lamdaOut => P(0)(801));
U_G1802: entity G port map(lamdaA => P(1)(290),lamdaB => P(1)(802),s => s(1)(290),lamdaOut => P(0)(802));
U_G1803: entity G port map(lamdaA => P(1)(291),lamdaB => P(1)(803),s => s(1)(291),lamdaOut => P(0)(803));
U_G1804: entity G port map(lamdaA => P(1)(292),lamdaB => P(1)(804),s => s(1)(292),lamdaOut => P(0)(804));
U_G1805: entity G port map(lamdaA => P(1)(293),lamdaB => P(1)(805),s => s(1)(293),lamdaOut => P(0)(805));
U_G1806: entity G port map(lamdaA => P(1)(294),lamdaB => P(1)(806),s => s(1)(294),lamdaOut => P(0)(806));
U_G1807: entity G port map(lamdaA => P(1)(295),lamdaB => P(1)(807),s => s(1)(295),lamdaOut => P(0)(807));
U_G1808: entity G port map(lamdaA => P(1)(296),lamdaB => P(1)(808),s => s(1)(296),lamdaOut => P(0)(808));
U_G1809: entity G port map(lamdaA => P(1)(297),lamdaB => P(1)(809),s => s(1)(297),lamdaOut => P(0)(809));
U_G1810: entity G port map(lamdaA => P(1)(298),lamdaB => P(1)(810),s => s(1)(298),lamdaOut => P(0)(810));
U_G1811: entity G port map(lamdaA => P(1)(299),lamdaB => P(1)(811),s => s(1)(299),lamdaOut => P(0)(811));
U_G1812: entity G port map(lamdaA => P(1)(300),lamdaB => P(1)(812),s => s(1)(300),lamdaOut => P(0)(812));
U_G1813: entity G port map(lamdaA => P(1)(301),lamdaB => P(1)(813),s => s(1)(301),lamdaOut => P(0)(813));
U_G1814: entity G port map(lamdaA => P(1)(302),lamdaB => P(1)(814),s => s(1)(302),lamdaOut => P(0)(814));
U_G1815: entity G port map(lamdaA => P(1)(303),lamdaB => P(1)(815),s => s(1)(303),lamdaOut => P(0)(815));
U_G1816: entity G port map(lamdaA => P(1)(304),lamdaB => P(1)(816),s => s(1)(304),lamdaOut => P(0)(816));
U_G1817: entity G port map(lamdaA => P(1)(305),lamdaB => P(1)(817),s => s(1)(305),lamdaOut => P(0)(817));
U_G1818: entity G port map(lamdaA => P(1)(306),lamdaB => P(1)(818),s => s(1)(306),lamdaOut => P(0)(818));
U_G1819: entity G port map(lamdaA => P(1)(307),lamdaB => P(1)(819),s => s(1)(307),lamdaOut => P(0)(819));
U_G1820: entity G port map(lamdaA => P(1)(308),lamdaB => P(1)(820),s => s(1)(308),lamdaOut => P(0)(820));
U_G1821: entity G port map(lamdaA => P(1)(309),lamdaB => P(1)(821),s => s(1)(309),lamdaOut => P(0)(821));
U_G1822: entity G port map(lamdaA => P(1)(310),lamdaB => P(1)(822),s => s(1)(310),lamdaOut => P(0)(822));
U_G1823: entity G port map(lamdaA => P(1)(311),lamdaB => P(1)(823),s => s(1)(311),lamdaOut => P(0)(823));
U_G1824: entity G port map(lamdaA => P(1)(312),lamdaB => P(1)(824),s => s(1)(312),lamdaOut => P(0)(824));
U_G1825: entity G port map(lamdaA => P(1)(313),lamdaB => P(1)(825),s => s(1)(313),lamdaOut => P(0)(825));
U_G1826: entity G port map(lamdaA => P(1)(314),lamdaB => P(1)(826),s => s(1)(314),lamdaOut => P(0)(826));
U_G1827: entity G port map(lamdaA => P(1)(315),lamdaB => P(1)(827),s => s(1)(315),lamdaOut => P(0)(827));
U_G1828: entity G port map(lamdaA => P(1)(316),lamdaB => P(1)(828),s => s(1)(316),lamdaOut => P(0)(828));
U_G1829: entity G port map(lamdaA => P(1)(317),lamdaB => P(1)(829),s => s(1)(317),lamdaOut => P(0)(829));
U_G1830: entity G port map(lamdaA => P(1)(318),lamdaB => P(1)(830),s => s(1)(318),lamdaOut => P(0)(830));
U_G1831: entity G port map(lamdaA => P(1)(319),lamdaB => P(1)(831),s => s(1)(319),lamdaOut => P(0)(831));
U_G1832: entity G port map(lamdaA => P(1)(320),lamdaB => P(1)(832),s => s(1)(320),lamdaOut => P(0)(832));
U_G1833: entity G port map(lamdaA => P(1)(321),lamdaB => P(1)(833),s => s(1)(321),lamdaOut => P(0)(833));
U_G1834: entity G port map(lamdaA => P(1)(322),lamdaB => P(1)(834),s => s(1)(322),lamdaOut => P(0)(834));
U_G1835: entity G port map(lamdaA => P(1)(323),lamdaB => P(1)(835),s => s(1)(323),lamdaOut => P(0)(835));
U_G1836: entity G port map(lamdaA => P(1)(324),lamdaB => P(1)(836),s => s(1)(324),lamdaOut => P(0)(836));
U_G1837: entity G port map(lamdaA => P(1)(325),lamdaB => P(1)(837),s => s(1)(325),lamdaOut => P(0)(837));
U_G1838: entity G port map(lamdaA => P(1)(326),lamdaB => P(1)(838),s => s(1)(326),lamdaOut => P(0)(838));
U_G1839: entity G port map(lamdaA => P(1)(327),lamdaB => P(1)(839),s => s(1)(327),lamdaOut => P(0)(839));
U_G1840: entity G port map(lamdaA => P(1)(328),lamdaB => P(1)(840),s => s(1)(328),lamdaOut => P(0)(840));
U_G1841: entity G port map(lamdaA => P(1)(329),lamdaB => P(1)(841),s => s(1)(329),lamdaOut => P(0)(841));
U_G1842: entity G port map(lamdaA => P(1)(330),lamdaB => P(1)(842),s => s(1)(330),lamdaOut => P(0)(842));
U_G1843: entity G port map(lamdaA => P(1)(331),lamdaB => P(1)(843),s => s(1)(331),lamdaOut => P(0)(843));
U_G1844: entity G port map(lamdaA => P(1)(332),lamdaB => P(1)(844),s => s(1)(332),lamdaOut => P(0)(844));
U_G1845: entity G port map(lamdaA => P(1)(333),lamdaB => P(1)(845),s => s(1)(333),lamdaOut => P(0)(845));
U_G1846: entity G port map(lamdaA => P(1)(334),lamdaB => P(1)(846),s => s(1)(334),lamdaOut => P(0)(846));
U_G1847: entity G port map(lamdaA => P(1)(335),lamdaB => P(1)(847),s => s(1)(335),lamdaOut => P(0)(847));
U_G1848: entity G port map(lamdaA => P(1)(336),lamdaB => P(1)(848),s => s(1)(336),lamdaOut => P(0)(848));
U_G1849: entity G port map(lamdaA => P(1)(337),lamdaB => P(1)(849),s => s(1)(337),lamdaOut => P(0)(849));
U_G1850: entity G port map(lamdaA => P(1)(338),lamdaB => P(1)(850),s => s(1)(338),lamdaOut => P(0)(850));
U_G1851: entity G port map(lamdaA => P(1)(339),lamdaB => P(1)(851),s => s(1)(339),lamdaOut => P(0)(851));
U_G1852: entity G port map(lamdaA => P(1)(340),lamdaB => P(1)(852),s => s(1)(340),lamdaOut => P(0)(852));
U_G1853: entity G port map(lamdaA => P(1)(341),lamdaB => P(1)(853),s => s(1)(341),lamdaOut => P(0)(853));
U_G1854: entity G port map(lamdaA => P(1)(342),lamdaB => P(1)(854),s => s(1)(342),lamdaOut => P(0)(854));
U_G1855: entity G port map(lamdaA => P(1)(343),lamdaB => P(1)(855),s => s(1)(343),lamdaOut => P(0)(855));
U_G1856: entity G port map(lamdaA => P(1)(344),lamdaB => P(1)(856),s => s(1)(344),lamdaOut => P(0)(856));
U_G1857: entity G port map(lamdaA => P(1)(345),lamdaB => P(1)(857),s => s(1)(345),lamdaOut => P(0)(857));
U_G1858: entity G port map(lamdaA => P(1)(346),lamdaB => P(1)(858),s => s(1)(346),lamdaOut => P(0)(858));
U_G1859: entity G port map(lamdaA => P(1)(347),lamdaB => P(1)(859),s => s(1)(347),lamdaOut => P(0)(859));
U_G1860: entity G port map(lamdaA => P(1)(348),lamdaB => P(1)(860),s => s(1)(348),lamdaOut => P(0)(860));
U_G1861: entity G port map(lamdaA => P(1)(349),lamdaB => P(1)(861),s => s(1)(349),lamdaOut => P(0)(861));
U_G1862: entity G port map(lamdaA => P(1)(350),lamdaB => P(1)(862),s => s(1)(350),lamdaOut => P(0)(862));
U_G1863: entity G port map(lamdaA => P(1)(351),lamdaB => P(1)(863),s => s(1)(351),lamdaOut => P(0)(863));
U_G1864: entity G port map(lamdaA => P(1)(352),lamdaB => P(1)(864),s => s(1)(352),lamdaOut => P(0)(864));
U_G1865: entity G port map(lamdaA => P(1)(353),lamdaB => P(1)(865),s => s(1)(353),lamdaOut => P(0)(865));
U_G1866: entity G port map(lamdaA => P(1)(354),lamdaB => P(1)(866),s => s(1)(354),lamdaOut => P(0)(866));
U_G1867: entity G port map(lamdaA => P(1)(355),lamdaB => P(1)(867),s => s(1)(355),lamdaOut => P(0)(867));
U_G1868: entity G port map(lamdaA => P(1)(356),lamdaB => P(1)(868),s => s(1)(356),lamdaOut => P(0)(868));
U_G1869: entity G port map(lamdaA => P(1)(357),lamdaB => P(1)(869),s => s(1)(357),lamdaOut => P(0)(869));
U_G1870: entity G port map(lamdaA => P(1)(358),lamdaB => P(1)(870),s => s(1)(358),lamdaOut => P(0)(870));
U_G1871: entity G port map(lamdaA => P(1)(359),lamdaB => P(1)(871),s => s(1)(359),lamdaOut => P(0)(871));
U_G1872: entity G port map(lamdaA => P(1)(360),lamdaB => P(1)(872),s => s(1)(360),lamdaOut => P(0)(872));
U_G1873: entity G port map(lamdaA => P(1)(361),lamdaB => P(1)(873),s => s(1)(361),lamdaOut => P(0)(873));
U_G1874: entity G port map(lamdaA => P(1)(362),lamdaB => P(1)(874),s => s(1)(362),lamdaOut => P(0)(874));
U_G1875: entity G port map(lamdaA => P(1)(363),lamdaB => P(1)(875),s => s(1)(363),lamdaOut => P(0)(875));
U_G1876: entity G port map(lamdaA => P(1)(364),lamdaB => P(1)(876),s => s(1)(364),lamdaOut => P(0)(876));
U_G1877: entity G port map(lamdaA => P(1)(365),lamdaB => P(1)(877),s => s(1)(365),lamdaOut => P(0)(877));
U_G1878: entity G port map(lamdaA => P(1)(366),lamdaB => P(1)(878),s => s(1)(366),lamdaOut => P(0)(878));
U_G1879: entity G port map(lamdaA => P(1)(367),lamdaB => P(1)(879),s => s(1)(367),lamdaOut => P(0)(879));
U_G1880: entity G port map(lamdaA => P(1)(368),lamdaB => P(1)(880),s => s(1)(368),lamdaOut => P(0)(880));
U_G1881: entity G port map(lamdaA => P(1)(369),lamdaB => P(1)(881),s => s(1)(369),lamdaOut => P(0)(881));
U_G1882: entity G port map(lamdaA => P(1)(370),lamdaB => P(1)(882),s => s(1)(370),lamdaOut => P(0)(882));
U_G1883: entity G port map(lamdaA => P(1)(371),lamdaB => P(1)(883),s => s(1)(371),lamdaOut => P(0)(883));
U_G1884: entity G port map(lamdaA => P(1)(372),lamdaB => P(1)(884),s => s(1)(372),lamdaOut => P(0)(884));
U_G1885: entity G port map(lamdaA => P(1)(373),lamdaB => P(1)(885),s => s(1)(373),lamdaOut => P(0)(885));
U_G1886: entity G port map(lamdaA => P(1)(374),lamdaB => P(1)(886),s => s(1)(374),lamdaOut => P(0)(886));
U_G1887: entity G port map(lamdaA => P(1)(375),lamdaB => P(1)(887),s => s(1)(375),lamdaOut => P(0)(887));
U_G1888: entity G port map(lamdaA => P(1)(376),lamdaB => P(1)(888),s => s(1)(376),lamdaOut => P(0)(888));
U_G1889: entity G port map(lamdaA => P(1)(377),lamdaB => P(1)(889),s => s(1)(377),lamdaOut => P(0)(889));
U_G1890: entity G port map(lamdaA => P(1)(378),lamdaB => P(1)(890),s => s(1)(378),lamdaOut => P(0)(890));
U_G1891: entity G port map(lamdaA => P(1)(379),lamdaB => P(1)(891),s => s(1)(379),lamdaOut => P(0)(891));
U_G1892: entity G port map(lamdaA => P(1)(380),lamdaB => P(1)(892),s => s(1)(380),lamdaOut => P(0)(892));
U_G1893: entity G port map(lamdaA => P(1)(381),lamdaB => P(1)(893),s => s(1)(381),lamdaOut => P(0)(893));
U_G1894: entity G port map(lamdaA => P(1)(382),lamdaB => P(1)(894),s => s(1)(382),lamdaOut => P(0)(894));
U_G1895: entity G port map(lamdaA => P(1)(383),lamdaB => P(1)(895),s => s(1)(383),lamdaOut => P(0)(895));
U_G1896: entity G port map(lamdaA => P(1)(384),lamdaB => P(1)(896),s => s(1)(384),lamdaOut => P(0)(896));
U_G1897: entity G port map(lamdaA => P(1)(385),lamdaB => P(1)(897),s => s(1)(385),lamdaOut => P(0)(897));
U_G1898: entity G port map(lamdaA => P(1)(386),lamdaB => P(1)(898),s => s(1)(386),lamdaOut => P(0)(898));
U_G1899: entity G port map(lamdaA => P(1)(387),lamdaB => P(1)(899),s => s(1)(387),lamdaOut => P(0)(899));
U_G1900: entity G port map(lamdaA => P(1)(388),lamdaB => P(1)(900),s => s(1)(388),lamdaOut => P(0)(900));
U_G1901: entity G port map(lamdaA => P(1)(389),lamdaB => P(1)(901),s => s(1)(389),lamdaOut => P(0)(901));
U_G1902: entity G port map(lamdaA => P(1)(390),lamdaB => P(1)(902),s => s(1)(390),lamdaOut => P(0)(902));
U_G1903: entity G port map(lamdaA => P(1)(391),lamdaB => P(1)(903),s => s(1)(391),lamdaOut => P(0)(903));
U_G1904: entity G port map(lamdaA => P(1)(392),lamdaB => P(1)(904),s => s(1)(392),lamdaOut => P(0)(904));
U_G1905: entity G port map(lamdaA => P(1)(393),lamdaB => P(1)(905),s => s(1)(393),lamdaOut => P(0)(905));
U_G1906: entity G port map(lamdaA => P(1)(394),lamdaB => P(1)(906),s => s(1)(394),lamdaOut => P(0)(906));
U_G1907: entity G port map(lamdaA => P(1)(395),lamdaB => P(1)(907),s => s(1)(395),lamdaOut => P(0)(907));
U_G1908: entity G port map(lamdaA => P(1)(396),lamdaB => P(1)(908),s => s(1)(396),lamdaOut => P(0)(908));
U_G1909: entity G port map(lamdaA => P(1)(397),lamdaB => P(1)(909),s => s(1)(397),lamdaOut => P(0)(909));
U_G1910: entity G port map(lamdaA => P(1)(398),lamdaB => P(1)(910),s => s(1)(398),lamdaOut => P(0)(910));
U_G1911: entity G port map(lamdaA => P(1)(399),lamdaB => P(1)(911),s => s(1)(399),lamdaOut => P(0)(911));
U_G1912: entity G port map(lamdaA => P(1)(400),lamdaB => P(1)(912),s => s(1)(400),lamdaOut => P(0)(912));
U_G1913: entity G port map(lamdaA => P(1)(401),lamdaB => P(1)(913),s => s(1)(401),lamdaOut => P(0)(913));
U_G1914: entity G port map(lamdaA => P(1)(402),lamdaB => P(1)(914),s => s(1)(402),lamdaOut => P(0)(914));
U_G1915: entity G port map(lamdaA => P(1)(403),lamdaB => P(1)(915),s => s(1)(403),lamdaOut => P(0)(915));
U_G1916: entity G port map(lamdaA => P(1)(404),lamdaB => P(1)(916),s => s(1)(404),lamdaOut => P(0)(916));
U_G1917: entity G port map(lamdaA => P(1)(405),lamdaB => P(1)(917),s => s(1)(405),lamdaOut => P(0)(917));
U_G1918: entity G port map(lamdaA => P(1)(406),lamdaB => P(1)(918),s => s(1)(406),lamdaOut => P(0)(918));
U_G1919: entity G port map(lamdaA => P(1)(407),lamdaB => P(1)(919),s => s(1)(407),lamdaOut => P(0)(919));
U_G1920: entity G port map(lamdaA => P(1)(408),lamdaB => P(1)(920),s => s(1)(408),lamdaOut => P(0)(920));
U_G1921: entity G port map(lamdaA => P(1)(409),lamdaB => P(1)(921),s => s(1)(409),lamdaOut => P(0)(921));
U_G1922: entity G port map(lamdaA => P(1)(410),lamdaB => P(1)(922),s => s(1)(410),lamdaOut => P(0)(922));
U_G1923: entity G port map(lamdaA => P(1)(411),lamdaB => P(1)(923),s => s(1)(411),lamdaOut => P(0)(923));
U_G1924: entity G port map(lamdaA => P(1)(412),lamdaB => P(1)(924),s => s(1)(412),lamdaOut => P(0)(924));
U_G1925: entity G port map(lamdaA => P(1)(413),lamdaB => P(1)(925),s => s(1)(413),lamdaOut => P(0)(925));
U_G1926: entity G port map(lamdaA => P(1)(414),lamdaB => P(1)(926),s => s(1)(414),lamdaOut => P(0)(926));
U_G1927: entity G port map(lamdaA => P(1)(415),lamdaB => P(1)(927),s => s(1)(415),lamdaOut => P(0)(927));
U_G1928: entity G port map(lamdaA => P(1)(416),lamdaB => P(1)(928),s => s(1)(416),lamdaOut => P(0)(928));
U_G1929: entity G port map(lamdaA => P(1)(417),lamdaB => P(1)(929),s => s(1)(417),lamdaOut => P(0)(929));
U_G1930: entity G port map(lamdaA => P(1)(418),lamdaB => P(1)(930),s => s(1)(418),lamdaOut => P(0)(930));
U_G1931: entity G port map(lamdaA => P(1)(419),lamdaB => P(1)(931),s => s(1)(419),lamdaOut => P(0)(931));
U_G1932: entity G port map(lamdaA => P(1)(420),lamdaB => P(1)(932),s => s(1)(420),lamdaOut => P(0)(932));
U_G1933: entity G port map(lamdaA => P(1)(421),lamdaB => P(1)(933),s => s(1)(421),lamdaOut => P(0)(933));
U_G1934: entity G port map(lamdaA => P(1)(422),lamdaB => P(1)(934),s => s(1)(422),lamdaOut => P(0)(934));
U_G1935: entity G port map(lamdaA => P(1)(423),lamdaB => P(1)(935),s => s(1)(423),lamdaOut => P(0)(935));
U_G1936: entity G port map(lamdaA => P(1)(424),lamdaB => P(1)(936),s => s(1)(424),lamdaOut => P(0)(936));
U_G1937: entity G port map(lamdaA => P(1)(425),lamdaB => P(1)(937),s => s(1)(425),lamdaOut => P(0)(937));
U_G1938: entity G port map(lamdaA => P(1)(426),lamdaB => P(1)(938),s => s(1)(426),lamdaOut => P(0)(938));
U_G1939: entity G port map(lamdaA => P(1)(427),lamdaB => P(1)(939),s => s(1)(427),lamdaOut => P(0)(939));
U_G1940: entity G port map(lamdaA => P(1)(428),lamdaB => P(1)(940),s => s(1)(428),lamdaOut => P(0)(940));
U_G1941: entity G port map(lamdaA => P(1)(429),lamdaB => P(1)(941),s => s(1)(429),lamdaOut => P(0)(941));
U_G1942: entity G port map(lamdaA => P(1)(430),lamdaB => P(1)(942),s => s(1)(430),lamdaOut => P(0)(942));
U_G1943: entity G port map(lamdaA => P(1)(431),lamdaB => P(1)(943),s => s(1)(431),lamdaOut => P(0)(943));
U_G1944: entity G port map(lamdaA => P(1)(432),lamdaB => P(1)(944),s => s(1)(432),lamdaOut => P(0)(944));
U_G1945: entity G port map(lamdaA => P(1)(433),lamdaB => P(1)(945),s => s(1)(433),lamdaOut => P(0)(945));
U_G1946: entity G port map(lamdaA => P(1)(434),lamdaB => P(1)(946),s => s(1)(434),lamdaOut => P(0)(946));
U_G1947: entity G port map(lamdaA => P(1)(435),lamdaB => P(1)(947),s => s(1)(435),lamdaOut => P(0)(947));
U_G1948: entity G port map(lamdaA => P(1)(436),lamdaB => P(1)(948),s => s(1)(436),lamdaOut => P(0)(948));
U_G1949: entity G port map(lamdaA => P(1)(437),lamdaB => P(1)(949),s => s(1)(437),lamdaOut => P(0)(949));
U_G1950: entity G port map(lamdaA => P(1)(438),lamdaB => P(1)(950),s => s(1)(438),lamdaOut => P(0)(950));
U_G1951: entity G port map(lamdaA => P(1)(439),lamdaB => P(1)(951),s => s(1)(439),lamdaOut => P(0)(951));
U_G1952: entity G port map(lamdaA => P(1)(440),lamdaB => P(1)(952),s => s(1)(440),lamdaOut => P(0)(952));
U_G1953: entity G port map(lamdaA => P(1)(441),lamdaB => P(1)(953),s => s(1)(441),lamdaOut => P(0)(953));
U_G1954: entity G port map(lamdaA => P(1)(442),lamdaB => P(1)(954),s => s(1)(442),lamdaOut => P(0)(954));
U_G1955: entity G port map(lamdaA => P(1)(443),lamdaB => P(1)(955),s => s(1)(443),lamdaOut => P(0)(955));
U_G1956: entity G port map(lamdaA => P(1)(444),lamdaB => P(1)(956),s => s(1)(444),lamdaOut => P(0)(956));
U_G1957: entity G port map(lamdaA => P(1)(445),lamdaB => P(1)(957),s => s(1)(445),lamdaOut => P(0)(957));
U_G1958: entity G port map(lamdaA => P(1)(446),lamdaB => P(1)(958),s => s(1)(446),lamdaOut => P(0)(958));
U_G1959: entity G port map(lamdaA => P(1)(447),lamdaB => P(1)(959),s => s(1)(447),lamdaOut => P(0)(959));
U_G1960: entity G port map(lamdaA => P(1)(448),lamdaB => P(1)(960),s => s(1)(448),lamdaOut => P(0)(960));
U_G1961: entity G port map(lamdaA => P(1)(449),lamdaB => P(1)(961),s => s(1)(449),lamdaOut => P(0)(961));
U_G1962: entity G port map(lamdaA => P(1)(450),lamdaB => P(1)(962),s => s(1)(450),lamdaOut => P(0)(962));
U_G1963: entity G port map(lamdaA => P(1)(451),lamdaB => P(1)(963),s => s(1)(451),lamdaOut => P(0)(963));
U_G1964: entity G port map(lamdaA => P(1)(452),lamdaB => P(1)(964),s => s(1)(452),lamdaOut => P(0)(964));
U_G1965: entity G port map(lamdaA => P(1)(453),lamdaB => P(1)(965),s => s(1)(453),lamdaOut => P(0)(965));
U_G1966: entity G port map(lamdaA => P(1)(454),lamdaB => P(1)(966),s => s(1)(454),lamdaOut => P(0)(966));
U_G1967: entity G port map(lamdaA => P(1)(455),lamdaB => P(1)(967),s => s(1)(455),lamdaOut => P(0)(967));
U_G1968: entity G port map(lamdaA => P(1)(456),lamdaB => P(1)(968),s => s(1)(456),lamdaOut => P(0)(968));
U_G1969: entity G port map(lamdaA => P(1)(457),lamdaB => P(1)(969),s => s(1)(457),lamdaOut => P(0)(969));
U_G1970: entity G port map(lamdaA => P(1)(458),lamdaB => P(1)(970),s => s(1)(458),lamdaOut => P(0)(970));
U_G1971: entity G port map(lamdaA => P(1)(459),lamdaB => P(1)(971),s => s(1)(459),lamdaOut => P(0)(971));
U_G1972: entity G port map(lamdaA => P(1)(460),lamdaB => P(1)(972),s => s(1)(460),lamdaOut => P(0)(972));
U_G1973: entity G port map(lamdaA => P(1)(461),lamdaB => P(1)(973),s => s(1)(461),lamdaOut => P(0)(973));
U_G1974: entity G port map(lamdaA => P(1)(462),lamdaB => P(1)(974),s => s(1)(462),lamdaOut => P(0)(974));
U_G1975: entity G port map(lamdaA => P(1)(463),lamdaB => P(1)(975),s => s(1)(463),lamdaOut => P(0)(975));
U_G1976: entity G port map(lamdaA => P(1)(464),lamdaB => P(1)(976),s => s(1)(464),lamdaOut => P(0)(976));
U_G1977: entity G port map(lamdaA => P(1)(465),lamdaB => P(1)(977),s => s(1)(465),lamdaOut => P(0)(977));
U_G1978: entity G port map(lamdaA => P(1)(466),lamdaB => P(1)(978),s => s(1)(466),lamdaOut => P(0)(978));
U_G1979: entity G port map(lamdaA => P(1)(467),lamdaB => P(1)(979),s => s(1)(467),lamdaOut => P(0)(979));
U_G1980: entity G port map(lamdaA => P(1)(468),lamdaB => P(1)(980),s => s(1)(468),lamdaOut => P(0)(980));
U_G1981: entity G port map(lamdaA => P(1)(469),lamdaB => P(1)(981),s => s(1)(469),lamdaOut => P(0)(981));
U_G1982: entity G port map(lamdaA => P(1)(470),lamdaB => P(1)(982),s => s(1)(470),lamdaOut => P(0)(982));
U_G1983: entity G port map(lamdaA => P(1)(471),lamdaB => P(1)(983),s => s(1)(471),lamdaOut => P(0)(983));
U_G1984: entity G port map(lamdaA => P(1)(472),lamdaB => P(1)(984),s => s(1)(472),lamdaOut => P(0)(984));
U_G1985: entity G port map(lamdaA => P(1)(473),lamdaB => P(1)(985),s => s(1)(473),lamdaOut => P(0)(985));
U_G1986: entity G port map(lamdaA => P(1)(474),lamdaB => P(1)(986),s => s(1)(474),lamdaOut => P(0)(986));
U_G1987: entity G port map(lamdaA => P(1)(475),lamdaB => P(1)(987),s => s(1)(475),lamdaOut => P(0)(987));
U_G1988: entity G port map(lamdaA => P(1)(476),lamdaB => P(1)(988),s => s(1)(476),lamdaOut => P(0)(988));
U_G1989: entity G port map(lamdaA => P(1)(477),lamdaB => P(1)(989),s => s(1)(477),lamdaOut => P(0)(989));
U_G1990: entity G port map(lamdaA => P(1)(478),lamdaB => P(1)(990),s => s(1)(478),lamdaOut => P(0)(990));
U_G1991: entity G port map(lamdaA => P(1)(479),lamdaB => P(1)(991),s => s(1)(479),lamdaOut => P(0)(991));
U_G1992: entity G port map(lamdaA => P(1)(480),lamdaB => P(1)(992),s => s(1)(480),lamdaOut => P(0)(992));
U_G1993: entity G port map(lamdaA => P(1)(481),lamdaB => P(1)(993),s => s(1)(481),lamdaOut => P(0)(993));
U_G1994: entity G port map(lamdaA => P(1)(482),lamdaB => P(1)(994),s => s(1)(482),lamdaOut => P(0)(994));
U_G1995: entity G port map(lamdaA => P(1)(483),lamdaB => P(1)(995),s => s(1)(483),lamdaOut => P(0)(995));
U_G1996: entity G port map(lamdaA => P(1)(484),lamdaB => P(1)(996),s => s(1)(484),lamdaOut => P(0)(996));
U_G1997: entity G port map(lamdaA => P(1)(485),lamdaB => P(1)(997),s => s(1)(485),lamdaOut => P(0)(997));
U_G1998: entity G port map(lamdaA => P(1)(486),lamdaB => P(1)(998),s => s(1)(486),lamdaOut => P(0)(998));
U_G1999: entity G port map(lamdaA => P(1)(487),lamdaB => P(1)(999),s => s(1)(487),lamdaOut => P(0)(999));
U_G11000: entity G port map(lamdaA => P(1)(488),lamdaB => P(1)(1000),s => s(1)(488),lamdaOut => P(0)(1000));
U_G11001: entity G port map(lamdaA => P(1)(489),lamdaB => P(1)(1001),s => s(1)(489),lamdaOut => P(0)(1001));
U_G11002: entity G port map(lamdaA => P(1)(490),lamdaB => P(1)(1002),s => s(1)(490),lamdaOut => P(0)(1002));
U_G11003: entity G port map(lamdaA => P(1)(491),lamdaB => P(1)(1003),s => s(1)(491),lamdaOut => P(0)(1003));
U_G11004: entity G port map(lamdaA => P(1)(492),lamdaB => P(1)(1004),s => s(1)(492),lamdaOut => P(0)(1004));
U_G11005: entity G port map(lamdaA => P(1)(493),lamdaB => P(1)(1005),s => s(1)(493),lamdaOut => P(0)(1005));
U_G11006: entity G port map(lamdaA => P(1)(494),lamdaB => P(1)(1006),s => s(1)(494),lamdaOut => P(0)(1006));
U_G11007: entity G port map(lamdaA => P(1)(495),lamdaB => P(1)(1007),s => s(1)(495),lamdaOut => P(0)(1007));
U_G11008: entity G port map(lamdaA => P(1)(496),lamdaB => P(1)(1008),s => s(1)(496),lamdaOut => P(0)(1008));
U_G11009: entity G port map(lamdaA => P(1)(497),lamdaB => P(1)(1009),s => s(1)(497),lamdaOut => P(0)(1009));
U_G11010: entity G port map(lamdaA => P(1)(498),lamdaB => P(1)(1010),s => s(1)(498),lamdaOut => P(0)(1010));
U_G11011: entity G port map(lamdaA => P(1)(499),lamdaB => P(1)(1011),s => s(1)(499),lamdaOut => P(0)(1011));
U_G11012: entity G port map(lamdaA => P(1)(500),lamdaB => P(1)(1012),s => s(1)(500),lamdaOut => P(0)(1012));
U_G11013: entity G port map(lamdaA => P(1)(501),lamdaB => P(1)(1013),s => s(1)(501),lamdaOut => P(0)(1013));
U_G11014: entity G port map(lamdaA => P(1)(502),lamdaB => P(1)(1014),s => s(1)(502),lamdaOut => P(0)(1014));
U_G11015: entity G port map(lamdaA => P(1)(503),lamdaB => P(1)(1015),s => s(1)(503),lamdaOut => P(0)(1015));
U_G11016: entity G port map(lamdaA => P(1)(504),lamdaB => P(1)(1016),s => s(1)(504),lamdaOut => P(0)(1016));
U_G11017: entity G port map(lamdaA => P(1)(505),lamdaB => P(1)(1017),s => s(1)(505),lamdaOut => P(0)(1017));
U_G11018: entity G port map(lamdaA => P(1)(506),lamdaB => P(1)(1018),s => s(1)(506),lamdaOut => P(0)(1018));
U_G11019: entity G port map(lamdaA => P(1)(507),lamdaB => P(1)(1019),s => s(1)(507),lamdaOut => P(0)(1019));
U_G11020: entity G port map(lamdaA => P(1)(508),lamdaB => P(1)(1020),s => s(1)(508),lamdaOut => P(0)(1020));
U_G11021: entity G port map(lamdaA => P(1)(509),lamdaB => P(1)(1021),s => s(1)(509),lamdaOut => P(0)(1021));
U_G11022: entity G port map(lamdaA => P(1)(510),lamdaB => P(1)(1022),s => s(1)(510),lamdaOut => P(0)(1022));
U_G11023: entity G port map(lamdaA => P(1)(511),lamdaB => P(1)(1023),s => s(1)(511),lamdaOut => P(0)(1023));
--Output Registers
ce_outputs <= '1';
U_D_FF0: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1012)(sign_bit),
q => outputs(0));

U_D_FF1: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1004)(sign_bit),
q => outputs(1));

U_D_FF2: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(476)(sign_bit),
q => outputs(2));

U_D_FF3: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(988)(sign_bit),
q => outputs(3));

U_D_FF4: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(828)(sign_bit),
q => outputs(4));

U_D_FF5: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(700)(sign_bit),
q => outputs(5));

U_D_FF6: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(444)(sign_bit),
q => outputs(6));

U_D_FF7: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(956)(sign_bit),
q => outputs(7));

U_D_FF8: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(636)(sign_bit),
q => outputs(8));

U_D_FF9: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(380)(sign_bit),
q => outputs(9));

U_D_FF10: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(892)(sign_bit),
q => outputs(10));

U_D_FF11: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(252)(sign_bit),
q => outputs(11));

U_D_FF12: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(764)(sign_bit),
q => outputs(12));

U_D_FF13: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(508)(sign_bit),
q => outputs(13));

U_D_FF14: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1020)(sign_bit),
q => outputs(14));

U_D_FF15: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1010)(sign_bit),
q => outputs(15));

U_D_FF16: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(874)(sign_bit),
q => outputs(16));

U_D_FF17: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(746)(sign_bit),
q => outputs(17));

U_D_FF18: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(490)(sign_bit),
q => outputs(18));

U_D_FF19: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1002)(sign_bit),
q => outputs(19));

U_D_FF20: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(922)(sign_bit),
q => outputs(20));

U_D_FF21: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(858)(sign_bit),
q => outputs(21));

U_D_FF22: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(730)(sign_bit),
q => outputs(22));

U_D_FF23: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(474)(sign_bit),
q => outputs(23));

U_D_FF24: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(986)(sign_bit),
q => outputs(24));

U_D_FF25: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(826)(sign_bit),
q => outputs(25));

U_D_FF26: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(186)(sign_bit),
q => outputs(26));

U_D_FF27: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(698)(sign_bit),
q => outputs(27));

U_D_FF28: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(442)(sign_bit),
q => outputs(28));

U_D_FF29: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(954)(sign_bit),
q => outputs(29));

U_D_FF30: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(122)(sign_bit),
q => outputs(30));

U_D_FF31: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(634)(sign_bit),
q => outputs(31));

U_D_FF32: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(378)(sign_bit),
q => outputs(32));

U_D_FF33: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(890)(sign_bit),
q => outputs(33));

U_D_FF34: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(250)(sign_bit),
q => outputs(34));

U_D_FF35: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(762)(sign_bit),
q => outputs(35));

U_D_FF36: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(506)(sign_bit),
q => outputs(36));

U_D_FF37: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1018)(sign_bit),
q => outputs(37));

U_D_FF38: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(966)(sign_bit),
q => outputs(38));

U_D_FF39: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(934)(sign_bit),
q => outputs(39));

U_D_FF40: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(870)(sign_bit),
q => outputs(40));

U_D_FF41: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(230)(sign_bit),
q => outputs(41));

U_D_FF42: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(742)(sign_bit),
q => outputs(42));

U_D_FF43: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(486)(sign_bit),
q => outputs(43));

U_D_FF44: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(998)(sign_bit),
q => outputs(44));

U_D_FF45: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(918)(sign_bit),
q => outputs(45));

U_D_FF46: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(598)(sign_bit),
q => outputs(46));

U_D_FF47: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(342)(sign_bit),
q => outputs(47));

U_D_FF48: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(854)(sign_bit),
q => outputs(48));

U_D_FF49: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(214)(sign_bit),
q => outputs(49));

U_D_FF50: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(726)(sign_bit),
q => outputs(50));

U_D_FF51: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(470)(sign_bit),
q => outputs(51));

U_D_FF52: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(982)(sign_bit),
q => outputs(52));

U_D_FF53: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(566)(sign_bit),
q => outputs(53));

U_D_FF54: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(310)(sign_bit),
q => outputs(54));

U_D_FF55: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(822)(sign_bit),
q => outputs(55));

U_D_FF56: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(182)(sign_bit),
q => outputs(56));

U_D_FF57: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(694)(sign_bit),
q => outputs(57));

U_D_FF58: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(438)(sign_bit),
q => outputs(58));

U_D_FF59: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(950)(sign_bit),
q => outputs(59));

U_D_FF60: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(118)(sign_bit),
q => outputs(60));

U_D_FF61: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(630)(sign_bit),
q => outputs(61));

U_D_FF62: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(374)(sign_bit),
q => outputs(62));

U_D_FF63: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(886)(sign_bit),
q => outputs(63));

U_D_FF64: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(246)(sign_bit),
q => outputs(64));

U_D_FF65: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(758)(sign_bit),
q => outputs(65));

U_D_FF66: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(502)(sign_bit),
q => outputs(66));

U_D_FF67: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1014)(sign_bit),
q => outputs(67));

U_D_FF68: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(782)(sign_bit),
q => outputs(68));

U_D_FF69: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(654)(sign_bit),
q => outputs(69));

U_D_FF70: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(398)(sign_bit),
q => outputs(70));

U_D_FF71: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(910)(sign_bit),
q => outputs(71));

U_D_FF72: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(590)(sign_bit),
q => outputs(72));

U_D_FF73: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(334)(sign_bit),
q => outputs(73));

U_D_FF74: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(846)(sign_bit),
q => outputs(74));

U_D_FF75: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(206)(sign_bit),
q => outputs(75));

U_D_FF76: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(718)(sign_bit),
q => outputs(76));

U_D_FF77: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(462)(sign_bit),
q => outputs(77));

U_D_FF78: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(974)(sign_bit),
q => outputs(78));

U_D_FF79: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(46)(sign_bit),
q => outputs(79));

U_D_FF80: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(558)(sign_bit),
q => outputs(80));

U_D_FF81: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(302)(sign_bit),
q => outputs(81));

U_D_FF82: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(814)(sign_bit),
q => outputs(82));

U_D_FF83: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(174)(sign_bit),
q => outputs(83));

U_D_FF84: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(686)(sign_bit),
q => outputs(84));

U_D_FF85: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(430)(sign_bit),
q => outputs(85));

U_D_FF86: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(942)(sign_bit),
q => outputs(86));

U_D_FF87: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(110)(sign_bit),
q => outputs(87));

U_D_FF88: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(622)(sign_bit),
q => outputs(88));

U_D_FF89: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(366)(sign_bit),
q => outputs(89));

U_D_FF90: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(878)(sign_bit),
q => outputs(90));

U_D_FF91: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(238)(sign_bit),
q => outputs(91));

U_D_FF92: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(750)(sign_bit),
q => outputs(92));

U_D_FF93: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(494)(sign_bit),
q => outputs(93));

U_D_FF94: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1006)(sign_bit),
q => outputs(94));

U_D_FF95: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(30)(sign_bit),
q => outputs(95));

U_D_FF96: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(542)(sign_bit),
q => outputs(96));

U_D_FF97: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(286)(sign_bit),
q => outputs(97));

U_D_FF98: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(798)(sign_bit),
q => outputs(98));

U_D_FF99: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(158)(sign_bit),
q => outputs(99));

U_D_FF100: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(670)(sign_bit),
q => outputs(100));

U_D_FF101: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(414)(sign_bit),
q => outputs(101));

U_D_FF102: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(926)(sign_bit),
q => outputs(102));

U_D_FF103: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(94)(sign_bit),
q => outputs(103));

U_D_FF104: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(606)(sign_bit),
q => outputs(104));

U_D_FF105: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(350)(sign_bit),
q => outputs(105));

U_D_FF106: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(862)(sign_bit),
q => outputs(106));

U_D_FF107: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(222)(sign_bit),
q => outputs(107));

U_D_FF108: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(734)(sign_bit),
q => outputs(108));

U_D_FF109: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(478)(sign_bit),
q => outputs(109));

U_D_FF110: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(990)(sign_bit),
q => outputs(110));

U_D_FF111: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(62)(sign_bit),
q => outputs(111));

U_D_FF112: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(574)(sign_bit),
q => outputs(112));

U_D_FF113: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(318)(sign_bit),
q => outputs(113));

U_D_FF114: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(830)(sign_bit),
q => outputs(114));

U_D_FF115: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(190)(sign_bit),
q => outputs(115));

U_D_FF116: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(702)(sign_bit),
q => outputs(116));

U_D_FF117: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(446)(sign_bit),
q => outputs(117));

U_D_FF118: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(958)(sign_bit),
q => outputs(118));

U_D_FF119: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(126)(sign_bit),
q => outputs(119));

U_D_FF120: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(638)(sign_bit),
q => outputs(120));

U_D_FF121: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(382)(sign_bit),
q => outputs(121));

U_D_FF122: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(894)(sign_bit),
q => outputs(122));

U_D_FF123: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(254)(sign_bit),
q => outputs(123));

U_D_FF124: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(766)(sign_bit),
q => outputs(124));

U_D_FF125: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(510)(sign_bit),
q => outputs(125));

U_D_FF126: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1022)(sign_bit),
q => outputs(126));

U_D_FF127: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(945)(sign_bit),
q => outputs(127));

U_D_FF128: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(881)(sign_bit),
q => outputs(128));

U_D_FF129: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(753)(sign_bit),
q => outputs(129));

U_D_FF130: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(497)(sign_bit),
q => outputs(130));

U_D_FF131: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1009)(sign_bit),
q => outputs(131));

U_D_FF132: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(969)(sign_bit),
q => outputs(132));

U_D_FF133: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(937)(sign_bit),
q => outputs(133));

U_D_FF134: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(617)(sign_bit),
q => outputs(134));

U_D_FF135: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(361)(sign_bit),
q => outputs(135));

U_D_FF136: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(873)(sign_bit),
q => outputs(136));

U_D_FF137: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(233)(sign_bit),
q => outputs(137));

U_D_FF138: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(745)(sign_bit),
q => outputs(138));

U_D_FF139: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(489)(sign_bit),
q => outputs(139));

U_D_FF140: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1001)(sign_bit),
q => outputs(140));

U_D_FF141: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(665)(sign_bit),
q => outputs(141));

U_D_FF142: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(409)(sign_bit),
q => outputs(142));

U_D_FF143: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(921)(sign_bit),
q => outputs(143));

U_D_FF144: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(601)(sign_bit),
q => outputs(144));

U_D_FF145: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(345)(sign_bit),
q => outputs(145));

U_D_FF146: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(857)(sign_bit),
q => outputs(146));

U_D_FF147: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(217)(sign_bit),
q => outputs(147));

U_D_FF148: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(729)(sign_bit),
q => outputs(148));

U_D_FF149: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(473)(sign_bit),
q => outputs(149));

U_D_FF150: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(985)(sign_bit),
q => outputs(150));

U_D_FF151: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(569)(sign_bit),
q => outputs(151));

U_D_FF152: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(313)(sign_bit),
q => outputs(152));

U_D_FF153: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(825)(sign_bit),
q => outputs(153));

U_D_FF154: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(185)(sign_bit),
q => outputs(154));

U_D_FF155: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(697)(sign_bit),
q => outputs(155));

U_D_FF156: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(441)(sign_bit),
q => outputs(156));

U_D_FF157: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(953)(sign_bit),
q => outputs(157));

U_D_FF158: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(121)(sign_bit),
q => outputs(158));

U_D_FF159: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(633)(sign_bit),
q => outputs(159));

U_D_FF160: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(377)(sign_bit),
q => outputs(160));

U_D_FF161: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(889)(sign_bit),
q => outputs(161));

U_D_FF162: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(249)(sign_bit),
q => outputs(162));

U_D_FF163: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(761)(sign_bit),
q => outputs(163));

U_D_FF164: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(505)(sign_bit),
q => outputs(164));

U_D_FF165: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1017)(sign_bit),
q => outputs(165));

U_D_FF166: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(709)(sign_bit),
q => outputs(166));

U_D_FF167: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(453)(sign_bit),
q => outputs(167));

U_D_FF168: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(965)(sign_bit),
q => outputs(168));

U_D_FF169: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(805)(sign_bit),
q => outputs(169));

U_D_FF170: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(677)(sign_bit),
q => outputs(170));

U_D_FF171: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(421)(sign_bit),
q => outputs(171));

U_D_FF172: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(933)(sign_bit),
q => outputs(172));

U_D_FF173: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(613)(sign_bit),
q => outputs(173));

U_D_FF174: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(357)(sign_bit),
q => outputs(174));

U_D_FF175: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(869)(sign_bit),
q => outputs(175));

U_D_FF176: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(229)(sign_bit),
q => outputs(176));

U_D_FF177: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(741)(sign_bit),
q => outputs(177));

U_D_FF178: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(485)(sign_bit),
q => outputs(178));

U_D_FF179: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(997)(sign_bit),
q => outputs(179));

U_D_FF180: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(789)(sign_bit),
q => outputs(180));

U_D_FF181: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(661)(sign_bit),
q => outputs(181));

U_D_FF182: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(405)(sign_bit),
q => outputs(182));

U_D_FF183: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(917)(sign_bit),
q => outputs(183));

U_D_FF184: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(85)(sign_bit),
q => outputs(184));

U_D_FF185: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(597)(sign_bit),
q => outputs(185));

U_D_FF186: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(341)(sign_bit),
q => outputs(186));

U_D_FF187: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(853)(sign_bit),
q => outputs(187));

U_D_FF188: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(213)(sign_bit),
q => outputs(188));

U_D_FF189: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(725)(sign_bit),
q => outputs(189));

U_D_FF190: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(469)(sign_bit),
q => outputs(190));

U_D_FF191: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(981)(sign_bit),
q => outputs(191));

U_D_FF192: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(53)(sign_bit),
q => outputs(192));

U_D_FF193: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(565)(sign_bit),
q => outputs(193));

U_D_FF194: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(309)(sign_bit),
q => outputs(194));

U_D_FF195: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(821)(sign_bit),
q => outputs(195));

U_D_FF196: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(181)(sign_bit),
q => outputs(196));

U_D_FF197: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(693)(sign_bit),
q => outputs(197));

U_D_FF198: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(437)(sign_bit),
q => outputs(198));

U_D_FF199: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(949)(sign_bit),
q => outputs(199));

U_D_FF200: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(117)(sign_bit),
q => outputs(200));

U_D_FF201: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(629)(sign_bit),
q => outputs(201));

U_D_FF202: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(373)(sign_bit),
q => outputs(202));

U_D_FF203: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(885)(sign_bit),
q => outputs(203));

U_D_FF204: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(245)(sign_bit),
q => outputs(204));

U_D_FF205: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(757)(sign_bit),
q => outputs(205));

U_D_FF206: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(501)(sign_bit),
q => outputs(206));

U_D_FF207: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1013)(sign_bit),
q => outputs(207));

U_D_FF208: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(525)(sign_bit),
q => outputs(208));

U_D_FF209: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(269)(sign_bit),
q => outputs(209));

U_D_FF210: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(781)(sign_bit),
q => outputs(210));

U_D_FF211: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(141)(sign_bit),
q => outputs(211));

U_D_FF212: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(653)(sign_bit),
q => outputs(212));

U_D_FF213: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(397)(sign_bit),
q => outputs(213));

U_D_FF214: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(909)(sign_bit),
q => outputs(214));

U_D_FF215: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(77)(sign_bit),
q => outputs(215));

U_D_FF216: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(589)(sign_bit),
q => outputs(216));

U_D_FF217: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(333)(sign_bit),
q => outputs(217));

U_D_FF218: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(845)(sign_bit),
q => outputs(218));

U_D_FF219: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(205)(sign_bit),
q => outputs(219));

U_D_FF220: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(717)(sign_bit),
q => outputs(220));

U_D_FF221: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(461)(sign_bit),
q => outputs(221));

U_D_FF222: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(973)(sign_bit),
q => outputs(222));

U_D_FF223: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(45)(sign_bit),
q => outputs(223));

U_D_FF224: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(557)(sign_bit),
q => outputs(224));

U_D_FF225: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(301)(sign_bit),
q => outputs(225));

U_D_FF226: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(813)(sign_bit),
q => outputs(226));

U_D_FF227: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(173)(sign_bit),
q => outputs(227));

U_D_FF228: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(685)(sign_bit),
q => outputs(228));

U_D_FF229: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(429)(sign_bit),
q => outputs(229));

U_D_FF230: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(941)(sign_bit),
q => outputs(230));

U_D_FF231: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(109)(sign_bit),
q => outputs(231));

U_D_FF232: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(621)(sign_bit),
q => outputs(232));

U_D_FF233: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(365)(sign_bit),
q => outputs(233));

U_D_FF234: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(877)(sign_bit),
q => outputs(234));

U_D_FF235: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(237)(sign_bit),
q => outputs(235));

U_D_FF236: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(749)(sign_bit),
q => outputs(236));

U_D_FF237: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(493)(sign_bit),
q => outputs(237));

U_D_FF238: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1005)(sign_bit),
q => outputs(238));

U_D_FF239: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(29)(sign_bit),
q => outputs(239));

U_D_FF240: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(541)(sign_bit),
q => outputs(240));

U_D_FF241: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(285)(sign_bit),
q => outputs(241));

U_D_FF242: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(797)(sign_bit),
q => outputs(242));

U_D_FF243: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(157)(sign_bit),
q => outputs(243));

U_D_FF244: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(669)(sign_bit),
q => outputs(244));

U_D_FF245: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(413)(sign_bit),
q => outputs(245));

U_D_FF246: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(925)(sign_bit),
q => outputs(246));

U_D_FF247: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(93)(sign_bit),
q => outputs(247));

U_D_FF248: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(605)(sign_bit),
q => outputs(248));

U_D_FF249: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(349)(sign_bit),
q => outputs(249));

U_D_FF250: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(861)(sign_bit),
q => outputs(250));

U_D_FF251: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(221)(sign_bit),
q => outputs(251));

U_D_FF252: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(733)(sign_bit),
q => outputs(252));

U_D_FF253: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(477)(sign_bit),
q => outputs(253));

U_D_FF254: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(989)(sign_bit),
q => outputs(254));

U_D_FF255: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(61)(sign_bit),
q => outputs(255));

U_D_FF256: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(573)(sign_bit),
q => outputs(256));

U_D_FF257: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(317)(sign_bit),
q => outputs(257));

U_D_FF258: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(829)(sign_bit),
q => outputs(258));

U_D_FF259: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(189)(sign_bit),
q => outputs(259));

U_D_FF260: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(701)(sign_bit),
q => outputs(260));

U_D_FF261: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(445)(sign_bit),
q => outputs(261));

U_D_FF262: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(957)(sign_bit),
q => outputs(262));

U_D_FF263: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(125)(sign_bit),
q => outputs(263));

U_D_FF264: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(637)(sign_bit),
q => outputs(264));

U_D_FF265: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(381)(sign_bit),
q => outputs(265));

U_D_FF266: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(893)(sign_bit),
q => outputs(266));

U_D_FF267: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(253)(sign_bit),
q => outputs(267));

U_D_FF268: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(765)(sign_bit),
q => outputs(268));

U_D_FF269: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(509)(sign_bit),
q => outputs(269));

U_D_FF270: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1021)(sign_bit),
q => outputs(270));

U_D_FF271: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(899)(sign_bit),
q => outputs(271));

U_D_FF272: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(835)(sign_bit),
q => outputs(272));

U_D_FF273: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(707)(sign_bit),
q => outputs(273));

U_D_FF274: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(451)(sign_bit),
q => outputs(274));

U_D_FF275: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(963)(sign_bit),
q => outputs(275));

U_D_FF276: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(291)(sign_bit),
q => outputs(276));

U_D_FF277: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(803)(sign_bit),
q => outputs(277));

U_D_FF278: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(163)(sign_bit),
q => outputs(278));

U_D_FF279: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(675)(sign_bit),
q => outputs(279));

U_D_FF280: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(419)(sign_bit),
q => outputs(280));

U_D_FF281: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(931)(sign_bit),
q => outputs(281));

U_D_FF282: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(99)(sign_bit),
q => outputs(282));

U_D_FF283: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(611)(sign_bit),
q => outputs(283));

U_D_FF284: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(355)(sign_bit),
q => outputs(284));

U_D_FF285: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(867)(sign_bit),
q => outputs(285));

U_D_FF286: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(227)(sign_bit),
q => outputs(286));

U_D_FF287: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(739)(sign_bit),
q => outputs(287));

U_D_FF288: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(483)(sign_bit),
q => outputs(288));

U_D_FF289: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(995)(sign_bit),
q => outputs(289));

U_D_FF290: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(531)(sign_bit),
q => outputs(290));

U_D_FF291: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(275)(sign_bit),
q => outputs(291));

U_D_FF292: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(787)(sign_bit),
q => outputs(292));

U_D_FF293: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(147)(sign_bit),
q => outputs(293));

U_D_FF294: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(659)(sign_bit),
q => outputs(294));

U_D_FF295: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(403)(sign_bit),
q => outputs(295));

U_D_FF296: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(915)(sign_bit),
q => outputs(296));

U_D_FF297: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(83)(sign_bit),
q => outputs(297));

U_D_FF298: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(595)(sign_bit),
q => outputs(298));

U_D_FF299: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(339)(sign_bit),
q => outputs(299));

U_D_FF300: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(851)(sign_bit),
q => outputs(300));

U_D_FF301: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(211)(sign_bit),
q => outputs(301));

U_D_FF302: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(723)(sign_bit),
q => outputs(302));

U_D_FF303: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(467)(sign_bit),
q => outputs(303));

U_D_FF304: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(979)(sign_bit),
q => outputs(304));

U_D_FF305: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(51)(sign_bit),
q => outputs(305));

U_D_FF306: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(563)(sign_bit),
q => outputs(306));

U_D_FF307: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(307)(sign_bit),
q => outputs(307));

U_D_FF308: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(819)(sign_bit),
q => outputs(308));

U_D_FF309: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(179)(sign_bit),
q => outputs(309));

U_D_FF310: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(691)(sign_bit),
q => outputs(310));

U_D_FF311: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(435)(sign_bit),
q => outputs(311));

U_D_FF312: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(947)(sign_bit),
q => outputs(312));

U_D_FF313: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(115)(sign_bit),
q => outputs(313));

U_D_FF314: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(627)(sign_bit),
q => outputs(314));

U_D_FF315: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(371)(sign_bit),
q => outputs(315));

U_D_FF316: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(883)(sign_bit),
q => outputs(316));

U_D_FF317: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(243)(sign_bit),
q => outputs(317));

U_D_FF318: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(755)(sign_bit),
q => outputs(318));

U_D_FF319: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(499)(sign_bit),
q => outputs(319));

U_D_FF320: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1011)(sign_bit),
q => outputs(320));

U_D_FF321: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(523)(sign_bit),
q => outputs(321));

U_D_FF322: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(267)(sign_bit),
q => outputs(322));

U_D_FF323: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(779)(sign_bit),
q => outputs(323));

U_D_FF324: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(139)(sign_bit),
q => outputs(324));

U_D_FF325: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(651)(sign_bit),
q => outputs(325));

U_D_FF326: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(395)(sign_bit),
q => outputs(326));

U_D_FF327: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(907)(sign_bit),
q => outputs(327));

U_D_FF328: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(75)(sign_bit),
q => outputs(328));

U_D_FF329: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(587)(sign_bit),
q => outputs(329));

U_D_FF330: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(331)(sign_bit),
q => outputs(330));

U_D_FF331: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(843)(sign_bit),
q => outputs(331));

U_D_FF332: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(203)(sign_bit),
q => outputs(332));

U_D_FF333: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(715)(sign_bit),
q => outputs(333));

U_D_FF334: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(459)(sign_bit),
q => outputs(334));

U_D_FF335: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(971)(sign_bit),
q => outputs(335));

U_D_FF336: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(43)(sign_bit),
q => outputs(336));

U_D_FF337: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(555)(sign_bit),
q => outputs(337));

U_D_FF338: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(299)(sign_bit),
q => outputs(338));

U_D_FF339: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(811)(sign_bit),
q => outputs(339));

U_D_FF340: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(171)(sign_bit),
q => outputs(340));

U_D_FF341: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(683)(sign_bit),
q => outputs(341));

U_D_FF342: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(427)(sign_bit),
q => outputs(342));

U_D_FF343: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(939)(sign_bit),
q => outputs(343));

U_D_FF344: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(107)(sign_bit),
q => outputs(344));

U_D_FF345: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(619)(sign_bit),
q => outputs(345));

U_D_FF346: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(363)(sign_bit),
q => outputs(346));

U_D_FF347: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(875)(sign_bit),
q => outputs(347));

U_D_FF348: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(235)(sign_bit),
q => outputs(348));

U_D_FF349: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(747)(sign_bit),
q => outputs(349));

U_D_FF350: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(491)(sign_bit),
q => outputs(350));

U_D_FF351: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1003)(sign_bit),
q => outputs(351));

U_D_FF352: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(27)(sign_bit),
q => outputs(352));

U_D_FF353: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(539)(sign_bit),
q => outputs(353));

U_D_FF354: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(283)(sign_bit),
q => outputs(354));

U_D_FF355: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(795)(sign_bit),
q => outputs(355));

U_D_FF356: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(155)(sign_bit),
q => outputs(356));

U_D_FF357: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(667)(sign_bit),
q => outputs(357));

U_D_FF358: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(411)(sign_bit),
q => outputs(358));

U_D_FF359: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(923)(sign_bit),
q => outputs(359));

U_D_FF360: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(91)(sign_bit),
q => outputs(360));

U_D_FF361: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(603)(sign_bit),
q => outputs(361));

U_D_FF362: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(347)(sign_bit),
q => outputs(362));

U_D_FF363: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(859)(sign_bit),
q => outputs(363));

U_D_FF364: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(219)(sign_bit),
q => outputs(364));

U_D_FF365: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(731)(sign_bit),
q => outputs(365));

U_D_FF366: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(475)(sign_bit),
q => outputs(366));

U_D_FF367: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(987)(sign_bit),
q => outputs(367));

U_D_FF368: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(59)(sign_bit),
q => outputs(368));

U_D_FF369: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(571)(sign_bit),
q => outputs(369));

U_D_FF370: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(315)(sign_bit),
q => outputs(370));

U_D_FF371: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(827)(sign_bit),
q => outputs(371));

U_D_FF372: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(187)(sign_bit),
q => outputs(372));

U_D_FF373: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(699)(sign_bit),
q => outputs(373));

U_D_FF374: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(443)(sign_bit),
q => outputs(374));

U_D_FF375: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(955)(sign_bit),
q => outputs(375));

U_D_FF376: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(123)(sign_bit),
q => outputs(376));

U_D_FF377: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(635)(sign_bit),
q => outputs(377));

U_D_FF378: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(379)(sign_bit),
q => outputs(378));

U_D_FF379: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(891)(sign_bit),
q => outputs(379));

U_D_FF380: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(251)(sign_bit),
q => outputs(380));

U_D_FF381: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(763)(sign_bit),
q => outputs(381));

U_D_FF382: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(507)(sign_bit),
q => outputs(382));

U_D_FF383: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1019)(sign_bit),
q => outputs(383));

U_D_FF384: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(7)(sign_bit),
q => outputs(384));

U_D_FF385: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(519)(sign_bit),
q => outputs(385));

U_D_FF386: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(263)(sign_bit),
q => outputs(386));

U_D_FF387: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(775)(sign_bit),
q => outputs(387));

U_D_FF388: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(135)(sign_bit),
q => outputs(388));

U_D_FF389: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(647)(sign_bit),
q => outputs(389));

U_D_FF390: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(391)(sign_bit),
q => outputs(390));

U_D_FF391: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(903)(sign_bit),
q => outputs(391));

U_D_FF392: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(71)(sign_bit),
q => outputs(392));

U_D_FF393: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(583)(sign_bit),
q => outputs(393));

U_D_FF394: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(327)(sign_bit),
q => outputs(394));

U_D_FF395: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(839)(sign_bit),
q => outputs(395));

U_D_FF396: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(199)(sign_bit),
q => outputs(396));

U_D_FF397: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(711)(sign_bit),
q => outputs(397));

U_D_FF398: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(455)(sign_bit),
q => outputs(398));

U_D_FF399: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(967)(sign_bit),
q => outputs(399));

U_D_FF400: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(39)(sign_bit),
q => outputs(400));

U_D_FF401: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(551)(sign_bit),
q => outputs(401));

U_D_FF402: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(295)(sign_bit),
q => outputs(402));

U_D_FF403: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(807)(sign_bit),
q => outputs(403));

U_D_FF404: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(167)(sign_bit),
q => outputs(404));

U_D_FF405: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(679)(sign_bit),
q => outputs(405));

U_D_FF406: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(423)(sign_bit),
q => outputs(406));

U_D_FF407: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(935)(sign_bit),
q => outputs(407));

U_D_FF408: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(103)(sign_bit),
q => outputs(408));

U_D_FF409: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(615)(sign_bit),
q => outputs(409));

U_D_FF410: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(359)(sign_bit),
q => outputs(410));

U_D_FF411: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(871)(sign_bit),
q => outputs(411));

U_D_FF412: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(231)(sign_bit),
q => outputs(412));

U_D_FF413: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(743)(sign_bit),
q => outputs(413));

U_D_FF414: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(487)(sign_bit),
q => outputs(414));

U_D_FF415: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(999)(sign_bit),
q => outputs(415));

U_D_FF416: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(23)(sign_bit),
q => outputs(416));

U_D_FF417: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(535)(sign_bit),
q => outputs(417));

U_D_FF418: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(279)(sign_bit),
q => outputs(418));

U_D_FF419: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(791)(sign_bit),
q => outputs(419));

U_D_FF420: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(151)(sign_bit),
q => outputs(420));

U_D_FF421: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(663)(sign_bit),
q => outputs(421));

U_D_FF422: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(407)(sign_bit),
q => outputs(422));

U_D_FF423: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(919)(sign_bit),
q => outputs(423));

U_D_FF424: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(87)(sign_bit),
q => outputs(424));

U_D_FF425: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(599)(sign_bit),
q => outputs(425));

U_D_FF426: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(343)(sign_bit),
q => outputs(426));

U_D_FF427: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(855)(sign_bit),
q => outputs(427));

U_D_FF428: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(215)(sign_bit),
q => outputs(428));

U_D_FF429: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(727)(sign_bit),
q => outputs(429));

U_D_FF430: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(471)(sign_bit),
q => outputs(430));

U_D_FF431: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(983)(sign_bit),
q => outputs(431));

U_D_FF432: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(55)(sign_bit),
q => outputs(432));

U_D_FF433: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(567)(sign_bit),
q => outputs(433));

U_D_FF434: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(311)(sign_bit),
q => outputs(434));

U_D_FF435: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(823)(sign_bit),
q => outputs(435));

U_D_FF436: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(183)(sign_bit),
q => outputs(436));

U_D_FF437: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(695)(sign_bit),
q => outputs(437));

U_D_FF438: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(439)(sign_bit),
q => outputs(438));

U_D_FF439: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(951)(sign_bit),
q => outputs(439));

U_D_FF440: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(119)(sign_bit),
q => outputs(440));

U_D_FF441: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(631)(sign_bit),
q => outputs(441));

U_D_FF442: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(375)(sign_bit),
q => outputs(442));

U_D_FF443: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(887)(sign_bit),
q => outputs(443));

U_D_FF444: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(247)(sign_bit),
q => outputs(444));

U_D_FF445: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(759)(sign_bit),
q => outputs(445));

U_D_FF446: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(503)(sign_bit),
q => outputs(446));

U_D_FF447: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1015)(sign_bit),
q => outputs(447));

U_D_FF448: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(15)(sign_bit),
q => outputs(448));

U_D_FF449: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(527)(sign_bit),
q => outputs(449));

U_D_FF450: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(271)(sign_bit),
q => outputs(450));

U_D_FF451: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(783)(sign_bit),
q => outputs(451));

U_D_FF452: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(143)(sign_bit),
q => outputs(452));

U_D_FF453: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(655)(sign_bit),
q => outputs(453));

U_D_FF454: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(399)(sign_bit),
q => outputs(454));

U_D_FF455: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(911)(sign_bit),
q => outputs(455));

U_D_FF456: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(79)(sign_bit),
q => outputs(456));

U_D_FF457: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(591)(sign_bit),
q => outputs(457));

U_D_FF458: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(335)(sign_bit),
q => outputs(458));

U_D_FF459: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(847)(sign_bit),
q => outputs(459));

U_D_FF460: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(207)(sign_bit),
q => outputs(460));

U_D_FF461: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(719)(sign_bit),
q => outputs(461));

U_D_FF462: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(463)(sign_bit),
q => outputs(462));

U_D_FF463: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(975)(sign_bit),
q => outputs(463));

U_D_FF464: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(47)(sign_bit),
q => outputs(464));

U_D_FF465: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(559)(sign_bit),
q => outputs(465));

U_D_FF466: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(303)(sign_bit),
q => outputs(466));

U_D_FF467: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(815)(sign_bit),
q => outputs(467));

U_D_FF468: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(175)(sign_bit),
q => outputs(468));

U_D_FF469: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(687)(sign_bit),
q => outputs(469));

U_D_FF470: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(431)(sign_bit),
q => outputs(470));

U_D_FF471: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(943)(sign_bit),
q => outputs(471));

U_D_FF472: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(111)(sign_bit),
q => outputs(472));

U_D_FF473: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(623)(sign_bit),
q => outputs(473));

U_D_FF474: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(367)(sign_bit),
q => outputs(474));

U_D_FF475: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(879)(sign_bit),
q => outputs(475));

U_D_FF476: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(239)(sign_bit),
q => outputs(476));

U_D_FF477: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(751)(sign_bit),
q => outputs(477));

U_D_FF478: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(495)(sign_bit),
q => outputs(478));

U_D_FF479: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1007)(sign_bit),
q => outputs(479));

U_D_FF480: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(31)(sign_bit),
q => outputs(480));

U_D_FF481: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(543)(sign_bit),
q => outputs(481));

U_D_FF482: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(287)(sign_bit),
q => outputs(482));

U_D_FF483: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(799)(sign_bit),
q => outputs(483));

U_D_FF484: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(159)(sign_bit),
q => outputs(484));

U_D_FF485: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(671)(sign_bit),
q => outputs(485));

U_D_FF486: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(415)(sign_bit),
q => outputs(486));

U_D_FF487: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(927)(sign_bit),
q => outputs(487));

U_D_FF488: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(95)(sign_bit),
q => outputs(488));

U_D_FF489: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(607)(sign_bit),
q => outputs(489));

U_D_FF490: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(351)(sign_bit),
q => outputs(490));

U_D_FF491: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(863)(sign_bit),
q => outputs(491));

U_D_FF492: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(223)(sign_bit),
q => outputs(492));

U_D_FF493: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(735)(sign_bit),
q => outputs(493));

U_D_FF494: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(479)(sign_bit),
q => outputs(494));

U_D_FF495: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(991)(sign_bit),
q => outputs(495));

U_D_FF496: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(63)(sign_bit),
q => outputs(496));

U_D_FF497: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(575)(sign_bit),
q => outputs(497));

U_D_FF498: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(319)(sign_bit),
q => outputs(498));

U_D_FF499: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(831)(sign_bit),
q => outputs(499));

U_D_FF500: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(191)(sign_bit),
q => outputs(500));

U_D_FF501: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(703)(sign_bit),
q => outputs(501));

U_D_FF502: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(447)(sign_bit),
q => outputs(502));

U_D_FF503: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(959)(sign_bit),
q => outputs(503));

U_D_FF504: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(127)(sign_bit),
q => outputs(504));

U_D_FF505: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(639)(sign_bit),
q => outputs(505));

U_D_FF506: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(383)(sign_bit),
q => outputs(506));

U_D_FF507: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(895)(sign_bit),
q => outputs(507));

U_D_FF508: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(255)(sign_bit),
q => outputs(508));

U_D_FF509: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(767)(sign_bit),
q => outputs(509));

U_D_FF510: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(511)(sign_bit),
q => outputs(510));

U_D_FF511: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(1023)(sign_bit),
q => outputs(511));
--Partial Sums Vector & Entity
u <=P(0)(511)(sign_bit)&P(0)(767)(sign_bit)&P(0)(255)(sign_bit)&P(0)(895)(sign_bit)&P(0)(383)(sign_bit)&P(0)(639)(sign_bit)&P(0)(127)(sign_bit)&P(0)(959)(sign_bit)&P(0)(447)(sign_bit)&P(0)(703)(sign_bit)&P(0)(191)(sign_bit)&P(0)(831)(sign_bit)&P(0)(319)(sign_bit)&P(0)(575)(sign_bit)&P(0)(63)(sign_bit)&P(0)(991)(sign_bit)&P(0)(479)(sign_bit)&P(0)(735)(sign_bit)&P(0)(223)(sign_bit)&P(0)(863)(sign_bit)&P(0)(351)(sign_bit)&P(0)(607)(sign_bit)&P(0)(95)(sign_bit)&P(0)(927)(sign_bit)&P(0)(415)(sign_bit)&P(0)(671)(sign_bit)&P(0)(159)(sign_bit)&P(0)(799)(sign_bit)&P(0)(287)(sign_bit)&P(0)(543)(sign_bit)&P(0)(31)(sign_bit)&P(0)(1007)(sign_bit)&P(0)(495)(sign_bit)&P(0)(751)(sign_bit)&P(0)(239)(sign_bit)&P(0)(879)(sign_bit)&P(0)(367)(sign_bit)&P(0)(623)(sign_bit)&P(0)(111)(sign_bit)&P(0)(943)(sign_bit)&P(0)(431)(sign_bit)&P(0)(687)(sign_bit)&P(0)(175)(sign_bit)&P(0)(815)(sign_bit)&P(0)(303)(sign_bit)&P(0)(559)(sign_bit)&P(0)(47)(sign_bit)&P(0)(975)(sign_bit)&P(0)(463)(sign_bit)&P(0)(719)(sign_bit)&P(0)(207)(sign_bit)&P(0)(847)(sign_bit)&P(0)(335)(sign_bit)&P(0)(591)(sign_bit)&P(0)(79)(sign_bit)&P(0)(911)(sign_bit)&P(0)(399)(sign_bit)&P(0)(655)(sign_bit)&P(0)(143)(sign_bit)&P(0)(783)(sign_bit)&P(0)(271)(sign_bit)&P(0)(527)(sign_bit)&P(0)(15)(sign_bit)&P(0)(1015)(sign_bit)&P(0)(503)(sign_bit)&P(0)(759)(sign_bit)&P(0)(247)(sign_bit)&P(0)(887)(sign_bit)&P(0)(375)(sign_bit)&P(0)(631)(sign_bit)&P(0)(119)(sign_bit)&P(0)(951)(sign_bit)&P(0)(439)(sign_bit)&P(0)(695)(sign_bit)&P(0)(183)(sign_bit)&P(0)(823)(sign_bit)&P(0)(311)(sign_bit)&P(0)(567)(sign_bit)&P(0)(55)(sign_bit)&P(0)(983)(sign_bit)&P(0)(471)(sign_bit)&P(0)(727)(sign_bit)&P(0)(215)(sign_bit)&P(0)(855)(sign_bit)&P(0)(343)(sign_bit)&P(0)(599)(sign_bit)&P(0)(87)(sign_bit)&P(0)(919)(sign_bit)&P(0)(407)(sign_bit)&P(0)(663)(sign_bit)&P(0)(151)(sign_bit)&P(0)(791)(sign_bit)&P(0)(279)(sign_bit)&P(0)(535)(sign_bit)&P(0)(23)(sign_bit)&P(0)(999)(sign_bit)&P(0)(487)(sign_bit)&P(0)(743)(sign_bit)&P(0)(231)(sign_bit)&P(0)(871)(sign_bit)&P(0)(359)(sign_bit)&P(0)(615)(sign_bit)&P(0)(103)(sign_bit)&P(0)(935)(sign_bit)&P(0)(423)(sign_bit)&P(0)(679)(sign_bit)&P(0)(167)(sign_bit)&P(0)(807)(sign_bit)&P(0)(295)(sign_bit)&P(0)(551)(sign_bit)&P(0)(39)(sign_bit)&P(0)(967)(sign_bit)&P(0)(455)(sign_bit)&P(0)(711)(sign_bit)&P(0)(199)(sign_bit)&P(0)(839)(sign_bit)&P(0)(327)(sign_bit)&P(0)(583)(sign_bit)&P(0)(71)(sign_bit)&P(0)(903)(sign_bit)&P(0)(391)(sign_bit)&P(0)(647)(sign_bit)&P(0)(135)(sign_bit)&P(0)(775)(sign_bit)&P(0)(263)(sign_bit)&P(0)(519)(sign_bit)&P(0)(7)(sign_bit)&P(0)(1019)(sign_bit)&P(0)(507)(sign_bit)&P(0)(763)(sign_bit)&P(0)(251)(sign_bit)&P(0)(891)(sign_bit)&P(0)(379)(sign_bit)&P(0)(635)(sign_bit)&P(0)(123)(sign_bit)&P(0)(955)(sign_bit)&P(0)(443)(sign_bit)&P(0)(699)(sign_bit)&P(0)(187)(sign_bit)&P(0)(827)(sign_bit)&P(0)(315)(sign_bit)&P(0)(571)(sign_bit)&P(0)(59)(sign_bit)&P(0)(987)(sign_bit)&P(0)(475)(sign_bit)&P(0)(731)(sign_bit)&P(0)(219)(sign_bit)&P(0)(859)(sign_bit)&P(0)(347)(sign_bit)&P(0)(603)(sign_bit)&P(0)(91)(sign_bit)&P(0)(923)(sign_bit)&P(0)(411)(sign_bit)&P(0)(667)(sign_bit)&P(0)(155)(sign_bit)&P(0)(795)(sign_bit)&P(0)(283)(sign_bit)&P(0)(539)(sign_bit)&P(0)(27)(sign_bit)&P(0)(1003)(sign_bit)&P(0)(491)(sign_bit)&P(0)(747)(sign_bit)&P(0)(235)(sign_bit)&P(0)(875)(sign_bit)&P(0)(363)(sign_bit)&P(0)(619)(sign_bit)&P(0)(107)(sign_bit)&P(0)(939)(sign_bit)&P(0)(427)(sign_bit)&P(0)(683)(sign_bit)&P(0)(171)(sign_bit)&P(0)(811)(sign_bit)&P(0)(299)(sign_bit)&P(0)(555)(sign_bit)&P(0)(43)(sign_bit)&P(0)(971)(sign_bit)&P(0)(459)(sign_bit)&P(0)(715)(sign_bit)&P(0)(203)(sign_bit)&P(0)(843)(sign_bit)&P(0)(331)(sign_bit)&P(0)(587)(sign_bit)&P(0)(75)(sign_bit)&P(0)(907)(sign_bit)&P(0)(395)(sign_bit)&P(0)(651)(sign_bit)&P(0)(139)(sign_bit)&P(0)(779)(sign_bit)&P(0)(267)(sign_bit)&P(0)(523)(sign_bit)&'0'&P(0)(1011)(sign_bit)&P(0)(499)(sign_bit)&P(0)(755)(sign_bit)&P(0)(243)(sign_bit)&P(0)(883)(sign_bit)&P(0)(371)(sign_bit)&P(0)(627)(sign_bit)&P(0)(115)(sign_bit)&P(0)(947)(sign_bit)&P(0)(435)(sign_bit)&P(0)(691)(sign_bit)&P(0)(179)(sign_bit)&P(0)(819)(sign_bit)&P(0)(307)(sign_bit)&P(0)(563)(sign_bit)&P(0)(51)(sign_bit)&P(0)(979)(sign_bit)&P(0)(467)(sign_bit)&P(0)(723)(sign_bit)&P(0)(211)(sign_bit)&P(0)(851)(sign_bit)&P(0)(339)(sign_bit)&P(0)(595)(sign_bit)&P(0)(83)(sign_bit)&P(0)(915)(sign_bit)&P(0)(403)(sign_bit)&P(0)(659)(sign_bit)&P(0)(147)(sign_bit)&P(0)(787)(sign_bit)&P(0)(275)(sign_bit)&P(0)(531)(sign_bit)&'0'&P(0)(995)(sign_bit)&P(0)(483)(sign_bit)&P(0)(739)(sign_bit)&P(0)(227)(sign_bit)&P(0)(867)(sign_bit)&P(0)(355)(sign_bit)&P(0)(611)(sign_bit)&P(0)(99)(sign_bit)&P(0)(931)(sign_bit)&P(0)(419)(sign_bit)&P(0)(675)(sign_bit)&P(0)(163)(sign_bit)&P(0)(803)(sign_bit)&P(0)(291)(sign_bit)&'0'&'0'&P(0)(963)(sign_bit)&P(0)(451)(sign_bit)&P(0)(707)(sign_bit)&'0'&P(0)(835)(sign_bit)&'0'&'0'&'0'&P(0)(899)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1021)(sign_bit)&P(0)(509)(sign_bit)&P(0)(765)(sign_bit)&P(0)(253)(sign_bit)&P(0)(893)(sign_bit)&P(0)(381)(sign_bit)&P(0)(637)(sign_bit)&P(0)(125)(sign_bit)&P(0)(957)(sign_bit)&P(0)(445)(sign_bit)&P(0)(701)(sign_bit)&P(0)(189)(sign_bit)&P(0)(829)(sign_bit)&P(0)(317)(sign_bit)&P(0)(573)(sign_bit)&P(0)(61)(sign_bit)&P(0)(989)(sign_bit)&P(0)(477)(sign_bit)&P(0)(733)(sign_bit)&P(0)(221)(sign_bit)&P(0)(861)(sign_bit)&P(0)(349)(sign_bit)&P(0)(605)(sign_bit)&P(0)(93)(sign_bit)&P(0)(925)(sign_bit)&P(0)(413)(sign_bit)&P(0)(669)(sign_bit)&P(0)(157)(sign_bit)&P(0)(797)(sign_bit)&P(0)(285)(sign_bit)&P(0)(541)(sign_bit)&P(0)(29)(sign_bit)&P(0)(1005)(sign_bit)&P(0)(493)(sign_bit)&P(0)(749)(sign_bit)&P(0)(237)(sign_bit)&P(0)(877)(sign_bit)&P(0)(365)(sign_bit)&P(0)(621)(sign_bit)&P(0)(109)(sign_bit)&P(0)(941)(sign_bit)&P(0)(429)(sign_bit)&P(0)(685)(sign_bit)&P(0)(173)(sign_bit)&P(0)(813)(sign_bit)&P(0)(301)(sign_bit)&P(0)(557)(sign_bit)&P(0)(45)(sign_bit)&P(0)(973)(sign_bit)&P(0)(461)(sign_bit)&P(0)(717)(sign_bit)&P(0)(205)(sign_bit)&P(0)(845)(sign_bit)&P(0)(333)(sign_bit)&P(0)(589)(sign_bit)&P(0)(77)(sign_bit)&P(0)(909)(sign_bit)&P(0)(397)(sign_bit)&P(0)(653)(sign_bit)&P(0)(141)(sign_bit)&P(0)(781)(sign_bit)&P(0)(269)(sign_bit)&P(0)(525)(sign_bit)&'0'&P(0)(1013)(sign_bit)&P(0)(501)(sign_bit)&P(0)(757)(sign_bit)&P(0)(245)(sign_bit)&P(0)(885)(sign_bit)&P(0)(373)(sign_bit)&P(0)(629)(sign_bit)&P(0)(117)(sign_bit)&P(0)(949)(sign_bit)&P(0)(437)(sign_bit)&P(0)(693)(sign_bit)&P(0)(181)(sign_bit)&P(0)(821)(sign_bit)&P(0)(309)(sign_bit)&P(0)(565)(sign_bit)&P(0)(53)(sign_bit)&P(0)(981)(sign_bit)&P(0)(469)(sign_bit)&P(0)(725)(sign_bit)&P(0)(213)(sign_bit)&P(0)(853)(sign_bit)&P(0)(341)(sign_bit)&P(0)(597)(sign_bit)&P(0)(85)(sign_bit)&P(0)(917)(sign_bit)&P(0)(405)(sign_bit)&P(0)(661)(sign_bit)&'0'&P(0)(789)(sign_bit)&'0'&'0'&'0'&P(0)(997)(sign_bit)&P(0)(485)(sign_bit)&P(0)(741)(sign_bit)&P(0)(229)(sign_bit)&P(0)(869)(sign_bit)&P(0)(357)(sign_bit)&P(0)(613)(sign_bit)&'0'&P(0)(933)(sign_bit)&P(0)(421)(sign_bit)&P(0)(677)(sign_bit)&'0'&P(0)(805)(sign_bit)&'0'&'0'&'0'&P(0)(965)(sign_bit)&P(0)(453)(sign_bit)&P(0)(709)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1017)(sign_bit)&P(0)(505)(sign_bit)&P(0)(761)(sign_bit)&P(0)(249)(sign_bit)&P(0)(889)(sign_bit)&P(0)(377)(sign_bit)&P(0)(633)(sign_bit)&P(0)(121)(sign_bit)&P(0)(953)(sign_bit)&P(0)(441)(sign_bit)&P(0)(697)(sign_bit)&P(0)(185)(sign_bit)&P(0)(825)(sign_bit)&P(0)(313)(sign_bit)&P(0)(569)(sign_bit)&'0'&P(0)(985)(sign_bit)&P(0)(473)(sign_bit)&P(0)(729)(sign_bit)&P(0)(217)(sign_bit)&P(0)(857)(sign_bit)&P(0)(345)(sign_bit)&P(0)(601)(sign_bit)&'0'&P(0)(921)(sign_bit)&P(0)(409)(sign_bit)&P(0)(665)(sign_bit)&'0'&'0'&'0'&'0'&'0'&P(0)(1001)(sign_bit)&P(0)(489)(sign_bit)&P(0)(745)(sign_bit)&P(0)(233)(sign_bit)&P(0)(873)(sign_bit)&P(0)(361)(sign_bit)&P(0)(617)(sign_bit)&'0'&P(0)(937)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(969)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1009)(sign_bit)&P(0)(497)(sign_bit)&P(0)(753)(sign_bit)&'0'&P(0)(881)(sign_bit)&'0'&'0'&'0'&P(0)(945)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1022)(sign_bit)&P(0)(510)(sign_bit)&P(0)(766)(sign_bit)&P(0)(254)(sign_bit)&P(0)(894)(sign_bit)&P(0)(382)(sign_bit)&P(0)(638)(sign_bit)&P(0)(126)(sign_bit)&P(0)(958)(sign_bit)&P(0)(446)(sign_bit)&P(0)(702)(sign_bit)&P(0)(190)(sign_bit)&P(0)(830)(sign_bit)&P(0)(318)(sign_bit)&P(0)(574)(sign_bit)&P(0)(62)(sign_bit)&P(0)(990)(sign_bit)&P(0)(478)(sign_bit)&P(0)(734)(sign_bit)&P(0)(222)(sign_bit)&P(0)(862)(sign_bit)&P(0)(350)(sign_bit)&P(0)(606)(sign_bit)&P(0)(94)(sign_bit)&P(0)(926)(sign_bit)&P(0)(414)(sign_bit)&P(0)(670)(sign_bit)&P(0)(158)(sign_bit)&P(0)(798)(sign_bit)&P(0)(286)(sign_bit)&P(0)(542)(sign_bit)&P(0)(30)(sign_bit)&P(0)(1006)(sign_bit)&P(0)(494)(sign_bit)&P(0)(750)(sign_bit)&P(0)(238)(sign_bit)&P(0)(878)(sign_bit)&P(0)(366)(sign_bit)&P(0)(622)(sign_bit)&P(0)(110)(sign_bit)&P(0)(942)(sign_bit)&P(0)(430)(sign_bit)&P(0)(686)(sign_bit)&P(0)(174)(sign_bit)&P(0)(814)(sign_bit)&P(0)(302)(sign_bit)&P(0)(558)(sign_bit)&P(0)(46)(sign_bit)&P(0)(974)(sign_bit)&P(0)(462)(sign_bit)&P(0)(718)(sign_bit)&P(0)(206)(sign_bit)&P(0)(846)(sign_bit)&P(0)(334)(sign_bit)&P(0)(590)(sign_bit)&'0'&P(0)(910)(sign_bit)&P(0)(398)(sign_bit)&P(0)(654)(sign_bit)&'0'&P(0)(782)(sign_bit)&'0'&'0'&'0'&P(0)(1014)(sign_bit)&P(0)(502)(sign_bit)&P(0)(758)(sign_bit)&P(0)(246)(sign_bit)&P(0)(886)(sign_bit)&P(0)(374)(sign_bit)&P(0)(630)(sign_bit)&P(0)(118)(sign_bit)&P(0)(950)(sign_bit)&P(0)(438)(sign_bit)&P(0)(694)(sign_bit)&P(0)(182)(sign_bit)&P(0)(822)(sign_bit)&P(0)(310)(sign_bit)&P(0)(566)(sign_bit)&'0'&P(0)(982)(sign_bit)&P(0)(470)(sign_bit)&P(0)(726)(sign_bit)&P(0)(214)(sign_bit)&P(0)(854)(sign_bit)&P(0)(342)(sign_bit)&P(0)(598)(sign_bit)&'0'&P(0)(918)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(998)(sign_bit)&P(0)(486)(sign_bit)&P(0)(742)(sign_bit)&P(0)(230)(sign_bit)&P(0)(870)(sign_bit)&'0'&'0'&'0'&P(0)(934)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(966)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1018)(sign_bit)&P(0)(506)(sign_bit)&P(0)(762)(sign_bit)&P(0)(250)(sign_bit)&P(0)(890)(sign_bit)&P(0)(378)(sign_bit)&P(0)(634)(sign_bit)&P(0)(122)(sign_bit)&P(0)(954)(sign_bit)&P(0)(442)(sign_bit)&P(0)(698)(sign_bit)&P(0)(186)(sign_bit)&P(0)(826)(sign_bit)&'0'&'0'&'0'&P(0)(986)(sign_bit)&P(0)(474)(sign_bit)&P(0)(730)(sign_bit)&'0'&P(0)(858)(sign_bit)&'0'&'0'&'0'&P(0)(922)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1002)(sign_bit)&P(0)(490)(sign_bit)&P(0)(746)(sign_bit)&'0'&P(0)(874)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1010)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1020)(sign_bit)&P(0)(508)(sign_bit)&P(0)(764)(sign_bit)&P(0)(252)(sign_bit)&P(0)(892)(sign_bit)&P(0)(380)(sign_bit)&P(0)(636)(sign_bit)&'0'&P(0)(956)(sign_bit)&P(0)(444)(sign_bit)&P(0)(700)(sign_bit)&'0'&P(0)(828)(sign_bit)&'0'&'0'&'0'&P(0)(988)(sign_bit)&P(0)(476)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1004)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(1012)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
U_Partials: entity work.PartialSumGenerator port map(u,s);
end Behavioral;


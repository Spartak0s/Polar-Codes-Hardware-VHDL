library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

entity synt4 is
port( 
	  address1	: in signed (5 downto 0);
	  stoixeio1	: out signed (80-1 downto 0)
);
end synt4;


architecture struct of synt4 is

    type rom_type is array (35 downto 0) of signed (79 downto 0);
    constant stoixeia : rom_type :=("11111111111111111111101000101100010101000001101111100000000000000000000000000000",
"11111111111111111111101000010101111010111111101010010000000000000000000000000000",
"11111111111111111111100111111110011110101100010011000000000000000000000000000000",
"11111111111111111111100111100101111010001111110110001000000000000000000000000000",
"11111111111111111111100111001100001000101000001011100000000000000000000000000000",
"11111111111111111111100110110001000010101100111101101000000000000000000000000000",
"11111111111111111111100110010100100001010101110110100000000000000000000000000000",
"11111111111111111111100101110110011100001001111110101000000000000000000000000000",
"11111111111111111111100101010110101001111010110010000000000000000000000000000000",
"11111111111111111111100100110100111111101110010101010000000000000000000000000000",
"11111111111111111111100100010001010001011010001010100000000000000000000000000000",
"11111111111111111111100011101011010001001000011100011000000000000000000000000000",
"11111111111111111111100011000010101110100010010001010000000000000000000000000000",
"11111111111111111111100010010111010111100101010111111000000000000000000000000000",
"11111111111111111111100001101000110110000011000010110000000000000000000000000000",
"11111111111111111111100000110110110000010101110100110000000000000000000000000000",
"11111111111111111111100000000000100111110110001000110000000000000000000000000000",
"11111111111111111111011111000101111000111010010010000000000000000000000000000000",
"11111111111111111111011110000101110111111010100001110000000000000000000000000000",
"11111111111111111111011100111111110000000000100101110000000000000000000000000000",
"11111111111111111111011011110010100000100110100011111000000000000000000000000000",
"11111111111111111111011010011100111000101111101000111000000000000000000000000000",
"11111111111111111111011000111101010101000001111001101000000000000000000000000000",
"11111111111111111111010111010001110101000111001110001000000000000000000000000000",
"11111111111111111111010101010111110110010000010011101000000000000000000000000000",
"11111111111111111111010011001100000101111001101100101000000000000000000000000000",
"11111111111111111111010000101010010000111010000001101000000000000000000000000000",
"11111111111111111111001101101100110000101010000011111000000000000000000000000000",
"11111111111111111111001010001011110100100011000010111000000000000000000000000000",
"11111111111111111111000101111000000001101010000111011000000000000000000000000000",
"11111111111111111110111111100101110110011110010000010000000000000000000000000000",
"11111111111111111110101000000000100110010110001100111000000000000000000000000000",
"11111111111111110101100111010111000010111101111010111000000000000000000000000000",
"00000000000111110111101101000011100101011000000100000110001001010000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000");

begin

stoixeio1<=stoixeia(to_integer((unsigned(address1))));
end struct;

----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:19:12 04/01/2016 
-- Design Name: 
-- Module Name:    Encoder1024 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.all;
use work.MyPackage.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Encoder1024 is
	Port ( inputs : in  STD_LOGIC_VECTOR (N/2-1 downto 0);
          outputs : out STD_LOGIC_VECTOR (N-1 downto 0));
end Encoder1024;

architecture Behavioral of Encoder1024 is

begin
outputs(0) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(1) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(2) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(271) xor inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(3) <= inputs(271) xor inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(4) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(5) <= inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(6) <= inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(7) <= inputs(384) xor inputs(385) xor inputs(386) xor inputs(387) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(8) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(9) <= inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(10) <= inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(11) <= inputs(321) xor inputs(322) xor inputs(323) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(12) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(13) <= inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(14) <= inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(15) <= inputs(448) xor inputs(449) xor inputs(450) xor inputs(451) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(16) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(17) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(18) <= inputs(15) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(19) <= inputs(290) xor inputs(291) xor inputs(292) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(20) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(21) <= inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(22) <= inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(23) <= inputs(416) xor inputs(417) xor inputs(418) xor inputs(419) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(24) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(25) <= inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(26) <= inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(27) <= inputs(352) xor inputs(353) xor inputs(354) xor inputs(355) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(28) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(29) <= inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(30) <= inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(31) <= inputs(480) xor inputs(481) xor inputs(482) xor inputs(483) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(32) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(33) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(34) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(35) <= inputs(276) xor inputs(277) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(36) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(37) <= inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(38) <= inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(39) <= inputs(400) xor inputs(401) xor inputs(402) xor inputs(403) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(40) <= inputs(1) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(41) <= inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(42) <= inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(43) <= inputs(336) xor inputs(337) xor inputs(338) xor inputs(339) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(44) <= inputs(1) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(45) <= inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(46) <= inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(47) <= inputs(464) xor inputs(465) xor inputs(466) xor inputs(467) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(48) <= inputs(0) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(49) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(50) <= inputs(15) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(51) <= inputs(305) xor inputs(306) xor inputs(307) xor inputs(308) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(52) <= inputs(0) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(53) <= inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(54) <= inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(55) <= inputs(432) xor inputs(433) xor inputs(434) xor inputs(435) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(56) <= inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(57) <= inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(58) <= inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(59) <= inputs(368) xor inputs(369) xor inputs(370) xor inputs(371) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(60) <= inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(61) <= inputs(255) xor inputs(256) xor inputs(257) xor inputs(258) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(62) <= inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(63) <= inputs(496) xor inputs(497) xor inputs(498) xor inputs(499) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(64) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(65) <= inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(66) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(67) <= inputs(272) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(68) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(69) <= inputs(166) xor inputs(167) xor inputs(168) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(70) <= inputs(38) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(71) <= inputs(392) xor inputs(393) xor inputs(394) xor inputs(395) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(72) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(73) <= inputs(132) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(74) <= inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(75) <= inputs(328) xor inputs(329) xor inputs(330) xor inputs(331) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(76) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(77) <= inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(78) <= inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(79) <= inputs(456) xor inputs(457) xor inputs(458) xor inputs(459) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(80) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(81) <= inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(82) <= inputs(15) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(83) <= inputs(297) xor inputs(298) xor inputs(299) xor inputs(300) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(84) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(85) <= inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(86) <= inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(87) <= inputs(424) xor inputs(425) xor inputs(426) xor inputs(427) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(88) <= inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(89) <= inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(90) <= inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(91) <= inputs(360) xor inputs(361) xor inputs(362) xor inputs(363) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(92) <= inputs(2) xor inputs(3) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(93) <= inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(94) <= inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(95) <= inputs(488) xor inputs(489) xor inputs(490) xor inputs(491) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(96) <= inputs(0) xor inputs(1) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(97) <= inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(98) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(99) <= inputs(282) xor inputs(283) xor inputs(284) xor inputs(285) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(100) <= inputs(0) xor inputs(1) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(101) <= inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(102) <= inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(103) <= inputs(408) xor inputs(409) xor inputs(410) xor inputs(411) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(104) <= inputs(1) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(105) <= inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(106) <= inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(107) <= inputs(344) xor inputs(345) xor inputs(346) xor inputs(347) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(108) <= inputs(1) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(109) <= inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(110) <= inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(111) <= inputs(472) xor inputs(473) xor inputs(474) xor inputs(475) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(112) <= inputs(0) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(113) <= inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(114) <= inputs(15) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(115) <= inputs(313) xor inputs(314) xor inputs(315) xor inputs(316) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(116) <= inputs(0) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(117) <= inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(118) <= inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(119) <= inputs(440) xor inputs(441) xor inputs(442) xor inputs(443) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(120) <= inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(121) <= inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(122) <= inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(123) <= inputs(376) xor inputs(377) xor inputs(378) xor inputs(379) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(124) <= inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(125) <= inputs(263) xor inputs(264) xor inputs(265) xor inputs(266) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(126) <= inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(127) <= inputs(504) xor inputs(505) xor inputs(506) xor inputs(507) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(128) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(129) <= inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(130) <= inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(271) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(131) <= inputs(271) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(132) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(133) <= inputs(166) xor inputs(167) xor inputs(168) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(134) <= inputs(38) xor inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(135) <= inputs(388) xor inputs(389) xor inputs(390) xor inputs(391) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(136) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(137) <= inputs(132) xor inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(138) <= inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(139) <= inputs(324) xor inputs(325) xor inputs(326) xor inputs(327) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(140) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(141) <= inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(142) <= inputs(69) xor inputs(70) xor inputs(71) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(143) <= inputs(452) xor inputs(453) xor inputs(454) xor inputs(455) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(144) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(145) <= inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(146) <= inputs(15) xor inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(147) <= inputs(293) xor inputs(294) xor inputs(295) xor inputs(296) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(148) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(149) <= inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(150) <= inputs(45) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(151) <= inputs(420) xor inputs(421) xor inputs(422) xor inputs(423) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(152) <= inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(153) <= inputs(141) xor inputs(142) xor inputs(143) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(154) <= inputs(20) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(155) <= inputs(356) xor inputs(357) xor inputs(358) xor inputs(359) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(156) <= inputs(2) xor inputs(3) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(157) <= inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(158) <= inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(159) <= inputs(484) xor inputs(485) xor inputs(486) xor inputs(487) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(160) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(161) <= inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(162) <= inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(163) <= inputs(278) xor inputs(279) xor inputs(280) xor inputs(281) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(164) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(165) <= inputs(170) xor inputs(171) xor inputs(172) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(166) <= inputs(39) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(167) <= inputs(404) xor inputs(405) xor inputs(406) xor inputs(407) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(168) <= inputs(1) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(169) <= inputs(133) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(170) <= inputs(17) xor inputs(18) xor inputs(19) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(171) <= inputs(340) xor inputs(341) xor inputs(342) xor inputs(343) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(172) <= inputs(1) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(173) <= inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(174) <= inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(175) <= inputs(468) xor inputs(469) xor inputs(470) xor inputs(471) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(176) <= inputs(0) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(177) <= inputs(127) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(178) <= inputs(15) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(179) <= inputs(309) xor inputs(310) xor inputs(311) xor inputs(312) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(180) <= inputs(0) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(181) <= inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(182) <= inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(183) <= inputs(436) xor inputs(437) xor inputs(438) xor inputs(439) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(184) <= inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(185) <= inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(186) <= inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(187) <= inputs(372) xor inputs(373) xor inputs(374) xor inputs(375) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(188) <= inputs(5) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(189) <= inputs(259) xor inputs(260) xor inputs(261) xor inputs(262) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(190) <= inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(191) <= inputs(500) xor inputs(501) xor inputs(502) xor inputs(503) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(192) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(193) <= inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(194) <= inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(273) xor inputs(274) xor inputs(275) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(195) <= inputs(273) xor inputs(274) xor inputs(275) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(196) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(197) <= inputs(166) xor inputs(167) xor inputs(168) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(198) <= inputs(38) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(199) <= inputs(396) xor inputs(397) xor inputs(398) xor inputs(399) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(200) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(201) <= inputs(132) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(202) <= inputs(17) xor inputs(18) xor inputs(19) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(203) <= inputs(332) xor inputs(333) xor inputs(334) xor inputs(335) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(204) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(205) <= inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(206) <= inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(207) <= inputs(460) xor inputs(461) xor inputs(462) xor inputs(463) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(208) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(209) <= inputs(129) xor inputs(130) xor inputs(131) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(210) <= inputs(15) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(211) <= inputs(301) xor inputs(302) xor inputs(303) xor inputs(304) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(212) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(213) <= inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(214) <= inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(215) <= inputs(428) xor inputs(429) xor inputs(430) xor inputs(431) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(216) <= inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(217) <= inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(218) <= inputs(22) xor inputs(23) xor inputs(24) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(219) <= inputs(364) xor inputs(365) xor inputs(366) xor inputs(367) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(220) <= inputs(2) xor inputs(3) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(221) <= inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(222) <= inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(223) <= inputs(492) xor inputs(493) xor inputs(494) xor inputs(495) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(224) <= inputs(0) xor inputs(1) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(225) <= inputs(129) xor inputs(130) xor inputs(131) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(226) <= inputs(15) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(227) <= inputs(286) xor inputs(287) xor inputs(288) xor inputs(289) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(228) <= inputs(0) xor inputs(1) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(229) <= inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(230) <= inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(231) <= inputs(412) xor inputs(413) xor inputs(414) xor inputs(415) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(232) <= inputs(1) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(233) <= inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(234) <= inputs(17) xor inputs(18) xor inputs(19) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(235) <= inputs(348) xor inputs(349) xor inputs(350) xor inputs(351) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(236) <= inputs(1) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(237) <= inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(238) <= inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(239) <= inputs(476) xor inputs(477) xor inputs(478) xor inputs(479) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(240) <= inputs(0) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(241) <= inputs(129) xor inputs(130) xor inputs(131) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(242) <= inputs(15) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(243) <= inputs(317) xor inputs(318) xor inputs(319) xor inputs(320) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(244) <= inputs(0) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(245) <= inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(246) <= inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(247) <= inputs(444) xor inputs(445) xor inputs(446) xor inputs(447) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(248) <= inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(249) <= inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(250) <= inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(251) <= inputs(380) xor inputs(381) xor inputs(382) xor inputs(383) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(252) <= inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(253) <= inputs(267) xor inputs(268) xor inputs(269) xor inputs(270) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(254) <= inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(255) <= inputs(508) xor inputs(509) xor inputs(510) xor inputs(511) ;
outputs(256) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(257) <= inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(258) <= inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(271) xor inputs(272) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(259) <= inputs(271) xor inputs(272) xor inputs(274) xor inputs(275) xor inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(260) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(261) <= inputs(167) xor inputs(168) xor inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(262) <= inputs(38) xor inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(263) <= inputs(386) xor inputs(387) xor inputs(390) xor inputs(391) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(264) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(265) <= inputs(132) xor inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(266) <= inputs(16) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(267) <= inputs(322) xor inputs(323) xor inputs(326) xor inputs(327) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(268) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(269) <= inputs(209) xor inputs(210) xor inputs(213) xor inputs(214) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(270) <= inputs(68) xor inputs(70) xor inputs(71) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(271) <= inputs(450) xor inputs(451) xor inputs(454) xor inputs(455) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(272) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(273) <= inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(274) <= inputs(15) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(275) <= inputs(291) xor inputs(292) xor inputs(295) xor inputs(296) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(276) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(277) <= inputs(180) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(278) <= inputs(45) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(279) <= inputs(418) xor inputs(419) xor inputs(422) xor inputs(423) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(280) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(281) <= inputs(142) xor inputs(143) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(282) <= inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(283) <= inputs(354) xor inputs(355) xor inputs(358) xor inputs(359) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(284) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(285) <= inputs(241) xor inputs(242) xor inputs(245) xor inputs(246) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(286) <= inputs(97) xor inputs(98) xor inputs(101) xor inputs(102) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(287) <= inputs(482) xor inputs(483) xor inputs(486) xor inputs(487) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(288) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(289) <= inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(290) <= inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(291) <= inputs(276) xor inputs(277) xor inputs(280) xor inputs(281) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(292) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(293) <= inputs(169) xor inputs(171) xor inputs(172) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(294) <= inputs(39) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(295) <= inputs(402) xor inputs(403) xor inputs(406) xor inputs(407) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(296) <= inputs(1) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(297) <= inputs(133) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(298) <= inputs(16) xor inputs(18) xor inputs(19) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(299) <= inputs(338) xor inputs(339) xor inputs(342) xor inputs(343) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(300) <= inputs(1) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(301) <= inputs(225) xor inputs(226) xor inputs(229) xor inputs(230) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(302) <= inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(303) <= inputs(466) xor inputs(467) xor inputs(470) xor inputs(471) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(304) <= inputs(0) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(305) <= inputs(127) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(306) <= inputs(15) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(307) <= inputs(307) xor inputs(308) xor inputs(311) xor inputs(312) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(308) <= inputs(0) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(309) <= inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(310) <= inputs(54) xor inputs(55) xor inputs(58) xor inputs(59) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(311) <= inputs(434) xor inputs(435) xor inputs(438) xor inputs(439) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(312) <= inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(313) <= inputs(152) xor inputs(153) xor inputs(156) xor inputs(157) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(314) <= inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(315) <= inputs(370) xor inputs(371) xor inputs(374) xor inputs(375) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(316) <= inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(317) <= inputs(257) xor inputs(258) xor inputs(261) xor inputs(262) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(318) <= inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(319) <= inputs(498) xor inputs(499) xor inputs(502) xor inputs(503) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(320) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(272) xor inputs(274) xor inputs(275) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(321) <= inputs(128) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(272) xor inputs(274) xor inputs(275) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(322) <= inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(272) xor inputs(274) xor inputs(275) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(323) <= inputs(272) xor inputs(274) xor inputs(275) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(324) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(167) xor inputs(168) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(325) <= inputs(167) xor inputs(168) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(326) <= inputs(38) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(327) <= inputs(394) xor inputs(395) xor inputs(398) xor inputs(399) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(328) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(329) <= inputs(132) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(330) <= inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(331) <= inputs(330) xor inputs(331) xor inputs(334) xor inputs(335) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(332) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(333) <= inputs(217) xor inputs(218) xor inputs(221) xor inputs(222) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(334) <= inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(335) <= inputs(458) xor inputs(459) xor inputs(462) xor inputs(463) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(336) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(337) <= inputs(128) xor inputs(130) xor inputs(131) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(338) <= inputs(15) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(339) <= inputs(299) xor inputs(300) xor inputs(303) xor inputs(304) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(340) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(341) <= inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(342) <= inputs(47) xor inputs(48) xor inputs(51) xor inputs(52) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(343) <= inputs(426) xor inputs(427) xor inputs(430) xor inputs(431) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(344) <= inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(345) <= inputs(145) xor inputs(146) xor inputs(149) xor inputs(150) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(346) <= inputs(21) xor inputs(23) xor inputs(24) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(347) <= inputs(362) xor inputs(363) xor inputs(366) xor inputs(367) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(348) <= inputs(2) xor inputs(3) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(349) <= inputs(249) xor inputs(250) xor inputs(253) xor inputs(254) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(350) <= inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(351) <= inputs(490) xor inputs(491) xor inputs(494) xor inputs(495) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(352) <= inputs(0) xor inputs(1) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(353) <= inputs(128) xor inputs(130) xor inputs(131) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(354) <= inputs(15) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(355) <= inputs(284) xor inputs(285) xor inputs(288) xor inputs(289) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(356) <= inputs(0) xor inputs(1) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(40) xor inputs(43) xor inputs(44) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(357) <= inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(358) <= inputs(40) xor inputs(43) xor inputs(44) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(359) <= inputs(410) xor inputs(411) xor inputs(414) xor inputs(415) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(360) <= inputs(1) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(361) <= inputs(135) xor inputs(136) xor inputs(139) xor inputs(140) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(362) <= inputs(16) xor inputs(18) xor inputs(19) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(363) <= inputs(346) xor inputs(347) xor inputs(350) xor inputs(351) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(364) <= inputs(1) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(365) <= inputs(233) xor inputs(234) xor inputs(237) xor inputs(238) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(366) <= inputs(89) xor inputs(90) xor inputs(93) xor inputs(94) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(367) <= inputs(474) xor inputs(475) xor inputs(478) xor inputs(479) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(368) <= inputs(0) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(131) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(369) <= inputs(128) xor inputs(130) xor inputs(131) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(370) <= inputs(15) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(371) <= inputs(315) xor inputs(316) xor inputs(319) xor inputs(320) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(372) <= inputs(0) xor inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(373) <= inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(374) <= inputs(62) xor inputs(63) xor inputs(66) xor inputs(67) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(375) <= inputs(442) xor inputs(443) xor inputs(446) xor inputs(447) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(376) <= inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(377) <= inputs(160) xor inputs(161) xor inputs(164) xor inputs(165) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(378) <= inputs(32) xor inputs(33) xor inputs(36) xor inputs(37) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(379) <= inputs(378) xor inputs(379) xor inputs(382) xor inputs(383) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(380) <= inputs(9) xor inputs(10) xor inputs(13) xor inputs(14) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(381) <= inputs(265) xor inputs(266) xor inputs(269) xor inputs(270) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(382) <= inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(383) <= inputs(506) xor inputs(507) xor inputs(510) xor inputs(511) ;
outputs(384) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(274) xor inputs(275) xor inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(385) <= inputs(127) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(271) xor inputs(274) xor inputs(275) xor inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(386) <= inputs(15) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(271) xor inputs(274) xor inputs(275) xor inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(387) <= inputs(271) xor inputs(274) xor inputs(275) xor inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(388) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(167) xor inputs(168) xor inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(389) <= inputs(167) xor inputs(168) xor inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(390) <= inputs(38) xor inputs(39) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(391) <= inputs(390) xor inputs(391) xor inputs(398) xor inputs(399) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(392) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(393) <= inputs(132) xor inputs(133) xor inputs(139) xor inputs(140) xor inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(394) <= inputs(18) xor inputs(19) xor inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(395) <= inputs(326) xor inputs(327) xor inputs(334) xor inputs(335) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(396) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(397) <= inputs(213) xor inputs(214) xor inputs(221) xor inputs(222) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(398) <= inputs(70) xor inputs(71) xor inputs(77) xor inputs(78) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(399) <= inputs(454) xor inputs(455) xor inputs(462) xor inputs(463) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(400) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(130) xor inputs(131) xor inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(401) <= inputs(127) xor inputs(130) xor inputs(131) xor inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(402) <= inputs(15) xor inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(403) <= inputs(295) xor inputs(296) xor inputs(303) xor inputs(304) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(404) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(405) <= inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(406) <= inputs(45) xor inputs(51) xor inputs(52) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(407) <= inputs(422) xor inputs(423) xor inputs(430) xor inputs(431) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(408) <= inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(409) <= inputs(142) xor inputs(143) xor inputs(149) xor inputs(150) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(410) <= inputs(20) xor inputs(23) xor inputs(24) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(411) <= inputs(358) xor inputs(359) xor inputs(366) xor inputs(367) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(412) <= inputs(2) xor inputs(3) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(413) <= inputs(245) xor inputs(246) xor inputs(253) xor inputs(254) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(414) <= inputs(101) xor inputs(102) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(415) <= inputs(486) xor inputs(487) xor inputs(494) xor inputs(495) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(416) <= inputs(0) xor inputs(1) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(18) xor inputs(19) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(43) xor inputs(44) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(139) xor inputs(140) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(417) <= inputs(127) xor inputs(130) xor inputs(131) xor inputs(133) xor inputs(139) xor inputs(140) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(418) <= inputs(15) xor inputs(18) xor inputs(19) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(39) xor inputs(43) xor inputs(44) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(419) <= inputs(280) xor inputs(281) xor inputs(288) xor inputs(289) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(420) <= inputs(0) xor inputs(1) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(39) xor inputs(43) xor inputs(44) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(421) <= inputs(171) xor inputs(172) xor inputs(178) xor inputs(179) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(422) <= inputs(39) xor inputs(43) xor inputs(44) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(423) <= inputs(406) xor inputs(407) xor inputs(414) xor inputs(415) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(424) <= inputs(1) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(18) xor inputs(19) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(139) xor inputs(140) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(425) <= inputs(133) xor inputs(139) xor inputs(140) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(426) <= inputs(18) xor inputs(19) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(427) <= inputs(342) xor inputs(343) xor inputs(350) xor inputs(351) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(428) <= inputs(1) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(429) <= inputs(229) xor inputs(230) xor inputs(237) xor inputs(238) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(430) <= inputs(85) xor inputs(86) xor inputs(93) xor inputs(94) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(431) <= inputs(470) xor inputs(471) xor inputs(478) xor inputs(479) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(432) <= inputs(0) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(130) xor inputs(131) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(433) <= inputs(127) xor inputs(130) xor inputs(131) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(434) <= inputs(15) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(435) <= inputs(311) xor inputs(312) xor inputs(319) xor inputs(320) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(436) <= inputs(0) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(437) <= inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(438) <= inputs(58) xor inputs(59) xor inputs(66) xor inputs(67) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(439) <= inputs(438) xor inputs(439) xor inputs(446) xor inputs(447) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(440) <= inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(441) <= inputs(156) xor inputs(157) xor inputs(164) xor inputs(165) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(442) <= inputs(28) xor inputs(29) xor inputs(36) xor inputs(37) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(443) <= inputs(374) xor inputs(375) xor inputs(382) xor inputs(383) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(444) <= inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(445) <= inputs(261) xor inputs(262) xor inputs(269) xor inputs(270) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(446) <= inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(447) <= inputs(502) xor inputs(503) xor inputs(510) xor inputs(511) ;
outputs(448) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(18) xor inputs(19) xor inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(139) xor inputs(140) xor inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(178) xor inputs(179) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(274) xor inputs(275) xor inputs(288) xor inputs(289) xor inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(449) <= inputs(130) xor inputs(131) xor inputs(132) xor inputs(139) xor inputs(140) xor inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(167) xor inputs(168) xor inputs(178) xor inputs(179) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(274) xor inputs(275) xor inputs(288) xor inputs(289) xor inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(450) <= inputs(15) xor inputs(18) xor inputs(19) xor inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(274) xor inputs(275) xor inputs(288) xor inputs(289) xor inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(451) <= inputs(274) xor inputs(275) xor inputs(288) xor inputs(289) xor inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(452) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(167) xor inputs(168) xor inputs(178) xor inputs(179) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(453) <= inputs(167) xor inputs(168) xor inputs(178) xor inputs(179) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(454) <= inputs(38) xor inputs(43) xor inputs(44) xor inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(455) <= inputs(398) xor inputs(399) xor inputs(414) xor inputs(415) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(456) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(18) xor inputs(19) xor inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(132) xor inputs(139) xor inputs(140) xor inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(457) <= inputs(132) xor inputs(139) xor inputs(140) xor inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(458) <= inputs(18) xor inputs(19) xor inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(459) <= inputs(334) xor inputs(335) xor inputs(350) xor inputs(351) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(460) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(461) <= inputs(221) xor inputs(222) xor inputs(237) xor inputs(238) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(462) <= inputs(77) xor inputs(78) xor inputs(93) xor inputs(94) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(463) <= inputs(462) xor inputs(463) xor inputs(478) xor inputs(479) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(464) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(130) xor inputs(131) xor inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(465) <= inputs(130) xor inputs(131) xor inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(466) <= inputs(15) xor inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(467) <= inputs(303) xor inputs(304) xor inputs(319) xor inputs(320) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(468) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(469) <= inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(470) <= inputs(51) xor inputs(52) xor inputs(66) xor inputs(67) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(471) <= inputs(430) xor inputs(431) xor inputs(446) xor inputs(447) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(472) <= inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(473) <= inputs(149) xor inputs(150) xor inputs(164) xor inputs(165) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(474) <= inputs(23) xor inputs(24) xor inputs(36) xor inputs(37) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(475) <= inputs(366) xor inputs(367) xor inputs(382) xor inputs(383) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(476) <= inputs(2) xor inputs(3) xor inputs(13) xor inputs(14) xor inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(477) <= inputs(253) xor inputs(254) xor inputs(269) xor inputs(270) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(478) <= inputs(109) xor inputs(110) xor inputs(125) xor inputs(126) xor inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(479) <= inputs(494) xor inputs(495) xor inputs(510) xor inputs(511) ;
outputs(480) <= inputs(0) xor inputs(1) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(18) xor inputs(19) xor inputs(36) xor inputs(37) xor inputs(43) xor inputs(44) xor inputs(66) xor inputs(67) xor inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(130) xor inputs(131) xor inputs(139) xor inputs(140) xor inputs(164) xor inputs(165) xor inputs(178) xor inputs(179) xor inputs(206) xor inputs(207) xor inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(288) xor inputs(289) xor inputs(319) xor inputs(320) xor inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(481) <= inputs(130) xor inputs(131) xor inputs(139) xor inputs(140) xor inputs(164) xor inputs(165) xor inputs(178) xor inputs(179) xor inputs(206) xor inputs(207) xor inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(288) xor inputs(289) xor inputs(319) xor inputs(320) xor inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(482) <= inputs(15) xor inputs(18) xor inputs(19) xor inputs(36) xor inputs(37) xor inputs(43) xor inputs(44) xor inputs(66) xor inputs(67) xor inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(288) xor inputs(289) xor inputs(319) xor inputs(320) xor inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(483) <= inputs(288) xor inputs(289) xor inputs(319) xor inputs(320) xor inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(484) <= inputs(0) xor inputs(1) xor inputs(13) xor inputs(14) xor inputs(43) xor inputs(44) xor inputs(66) xor inputs(67) xor inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(178) xor inputs(179) xor inputs(206) xor inputs(207) xor inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(485) <= inputs(178) xor inputs(179) xor inputs(206) xor inputs(207) xor inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(486) <= inputs(43) xor inputs(44) xor inputs(66) xor inputs(67) xor inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(487) <= inputs(414) xor inputs(415) xor inputs(446) xor inputs(447) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(488) <= inputs(1) xor inputs(13) xor inputs(14) xor inputs(18) xor inputs(19) xor inputs(36) xor inputs(37) xor inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(139) xor inputs(140) xor inputs(164) xor inputs(165) xor inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(489) <= inputs(139) xor inputs(140) xor inputs(164) xor inputs(165) xor inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(490) <= inputs(18) xor inputs(19) xor inputs(36) xor inputs(37) xor inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(491) <= inputs(350) xor inputs(351) xor inputs(382) xor inputs(383) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(492) <= inputs(1) xor inputs(13) xor inputs(14) xor inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(493) <= inputs(237) xor inputs(238) xor inputs(269) xor inputs(270) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(494) <= inputs(93) xor inputs(94) xor inputs(125) xor inputs(126) xor inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(495) <= inputs(478) xor inputs(479) xor inputs(510) xor inputs(511) ;
outputs(496) <= inputs(0) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(36) xor inputs(37) xor inputs(66) xor inputs(67) xor inputs(125) xor inputs(126) xor inputs(130) xor inputs(131) xor inputs(164) xor inputs(165) xor inputs(206) xor inputs(207) xor inputs(269) xor inputs(270) xor inputs(319) xor inputs(320) xor inputs(382) xor inputs(383) xor inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(497) <= inputs(130) xor inputs(131) xor inputs(164) xor inputs(165) xor inputs(206) xor inputs(207) xor inputs(269) xor inputs(270) xor inputs(319) xor inputs(320) xor inputs(382) xor inputs(383) xor inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(498) <= inputs(15) xor inputs(36) xor inputs(37) xor inputs(66) xor inputs(67) xor inputs(125) xor inputs(126) xor inputs(319) xor inputs(320) xor inputs(382) xor inputs(383) xor inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(499) <= inputs(319) xor inputs(320) xor inputs(382) xor inputs(383) xor inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(500) <= inputs(0) xor inputs(13) xor inputs(14) xor inputs(66) xor inputs(67) xor inputs(125) xor inputs(126) xor inputs(206) xor inputs(207) xor inputs(269) xor inputs(270) xor inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(501) <= inputs(206) xor inputs(207) xor inputs(269) xor inputs(270) xor inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(502) <= inputs(66) xor inputs(67) xor inputs(125) xor inputs(126) xor inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(503) <= inputs(446) xor inputs(447) xor inputs(510) xor inputs(511) ;
outputs(504) <= inputs(13) xor inputs(14) xor inputs(36) xor inputs(37) xor inputs(125) xor inputs(126) xor inputs(164) xor inputs(165) xor inputs(269) xor inputs(270) xor inputs(382) xor inputs(383) xor inputs(510) xor inputs(511) ;
outputs(505) <= inputs(164) xor inputs(165) xor inputs(269) xor inputs(270) xor inputs(382) xor inputs(383) xor inputs(510) xor inputs(511) ;
outputs(506) <= inputs(36) xor inputs(37) xor inputs(125) xor inputs(126) xor inputs(382) xor inputs(383) xor inputs(510) xor inputs(511) ;
outputs(507) <= inputs(382) xor inputs(383) xor inputs(510) xor inputs(511) ;
outputs(508) <= inputs(13) xor inputs(14) xor inputs(125) xor inputs(126) xor inputs(269) xor inputs(270) xor inputs(510) xor inputs(511) ;
outputs(509) <= inputs(269) xor inputs(270) xor inputs(510) xor inputs(511) ;
outputs(510) <= inputs(125) xor inputs(126) xor inputs(510) xor inputs(511) ;
outputs(511) <= inputs(510) xor inputs(511) ;
outputs(512) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(273) xor inputs(275) xor inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(513) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(273) xor inputs(275) xor inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(514) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(271) xor inputs(272) xor inputs(273) xor inputs(275) xor inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(515) <= inputs(271) xor inputs(272) xor inputs(273) xor inputs(275) xor inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(516) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(166) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(517) <= inputs(166) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(518) <= inputs(38) xor inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(519) <= inputs(385) xor inputs(387) xor inputs(389) xor inputs(391) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(520) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(521) <= inputs(132) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(522) <= inputs(16) xor inputs(17) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(523) <= inputs(321) xor inputs(323) xor inputs(325) xor inputs(327) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(524) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(525) <= inputs(208) xor inputs(210) xor inputs(212) xor inputs(214) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(526) <= inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(527) <= inputs(449) xor inputs(451) xor inputs(453) xor inputs(455) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(528) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(529) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(530) <= inputs(15) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(531) <= inputs(290) xor inputs(292) xor inputs(294) xor inputs(296) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(532) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(533) <= inputs(180) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(534) <= inputs(45) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(535) <= inputs(417) xor inputs(419) xor inputs(421) xor inputs(423) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(536) <= inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(537) <= inputs(141) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(538) <= inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(539) <= inputs(353) xor inputs(355) xor inputs(357) xor inputs(359) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(540) <= inputs(3) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(541) <= inputs(240) xor inputs(242) xor inputs(244) xor inputs(246) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(542) <= inputs(96) xor inputs(98) xor inputs(100) xor inputs(102) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(543) <= inputs(481) xor inputs(483) xor inputs(485) xor inputs(487) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(544) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(545) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(546) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(547) <= inputs(277) xor inputs(279) xor inputs(281) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(548) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(549) <= inputs(169) xor inputs(170) xor inputs(172) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(550) <= inputs(39) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(551) <= inputs(401) xor inputs(403) xor inputs(405) xor inputs(407) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(552) <= inputs(1) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(553) <= inputs(133) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(554) <= inputs(16) xor inputs(17) xor inputs(19) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(555) <= inputs(337) xor inputs(339) xor inputs(341) xor inputs(343) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(556) <= inputs(1) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(557) <= inputs(224) xor inputs(226) xor inputs(228) xor inputs(230) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(558) <= inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(559) <= inputs(465) xor inputs(467) xor inputs(469) xor inputs(471) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(560) <= inputs(0) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(561) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(562) <= inputs(15) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(563) <= inputs(306) xor inputs(308) xor inputs(310) xor inputs(312) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(564) <= inputs(0) xor inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(565) <= inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(566) <= inputs(53) xor inputs(55) xor inputs(57) xor inputs(59) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(567) <= inputs(433) xor inputs(435) xor inputs(437) xor inputs(439) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(568) <= inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(569) <= inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(570) <= inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(571) <= inputs(369) xor inputs(371) xor inputs(373) xor inputs(375) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(572) <= inputs(4) xor inputs(5) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(573) <= inputs(256) xor inputs(258) xor inputs(260) xor inputs(262) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(574) <= inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(575) <= inputs(497) xor inputs(499) xor inputs(501) xor inputs(503) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(576) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(132) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(272) xor inputs(273) xor inputs(275) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(577) <= inputs(128) xor inputs(129) xor inputs(131) xor inputs(132) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(272) xor inputs(273) xor inputs(275) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(578) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(272) xor inputs(273) xor inputs(275) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(579) <= inputs(272) xor inputs(273) xor inputs(275) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(580) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(166) xor inputs(168) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(581) <= inputs(166) xor inputs(168) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(582) <= inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(583) <= inputs(393) xor inputs(395) xor inputs(397) xor inputs(399) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(584) <= inputs(1) xor inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(585) <= inputs(132) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(586) <= inputs(16) xor inputs(17) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(587) <= inputs(329) xor inputs(331) xor inputs(333) xor inputs(335) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(588) <= inputs(1) xor inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(589) <= inputs(216) xor inputs(218) xor inputs(220) xor inputs(222) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(590) <= inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(591) <= inputs(457) xor inputs(459) xor inputs(461) xor inputs(463) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(592) <= inputs(0) xor inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(593) <= inputs(128) xor inputs(129) xor inputs(131) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(594) <= inputs(15) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(595) <= inputs(298) xor inputs(300) xor inputs(302) xor inputs(304) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(596) <= inputs(0) xor inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(597) <= inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(598) <= inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(599) <= inputs(425) xor inputs(427) xor inputs(429) xor inputs(431) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(600) <= inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(601) <= inputs(144) xor inputs(146) xor inputs(148) xor inputs(150) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(602) <= inputs(21) xor inputs(22) xor inputs(24) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(603) <= inputs(361) xor inputs(363) xor inputs(365) xor inputs(367) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(604) <= inputs(3) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(605) <= inputs(248) xor inputs(250) xor inputs(252) xor inputs(254) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(606) <= inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(607) <= inputs(489) xor inputs(491) xor inputs(493) xor inputs(495) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(608) <= inputs(0) xor inputs(1) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(609) <= inputs(128) xor inputs(129) xor inputs(131) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(610) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(611) <= inputs(283) xor inputs(285) xor inputs(287) xor inputs(289) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(612) <= inputs(0) xor inputs(1) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(613) <= inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(614) <= inputs(40) xor inputs(42) xor inputs(44) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(615) <= inputs(409) xor inputs(411) xor inputs(413) xor inputs(415) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(616) <= inputs(1) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(17) xor inputs(19) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(617) <= inputs(134) xor inputs(136) xor inputs(138) xor inputs(140) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(618) <= inputs(16) xor inputs(17) xor inputs(19) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(619) <= inputs(345) xor inputs(347) xor inputs(349) xor inputs(351) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(620) <= inputs(1) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(621) <= inputs(232) xor inputs(234) xor inputs(236) xor inputs(238) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(622) <= inputs(88) xor inputs(90) xor inputs(92) xor inputs(94) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(623) <= inputs(473) xor inputs(475) xor inputs(477) xor inputs(479) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(624) <= inputs(0) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(129) xor inputs(131) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(625) <= inputs(128) xor inputs(129) xor inputs(131) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(626) <= inputs(15) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(627) <= inputs(314) xor inputs(316) xor inputs(318) xor inputs(320) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(628) <= inputs(0) xor inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(629) <= inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(630) <= inputs(61) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(631) <= inputs(441) xor inputs(443) xor inputs(445) xor inputs(447) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(632) <= inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(633) <= inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(634) <= inputs(31) xor inputs(33) xor inputs(35) xor inputs(37) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(635) <= inputs(377) xor inputs(379) xor inputs(381) xor inputs(383) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(636) <= inputs(8) xor inputs(10) xor inputs(12) xor inputs(14) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(637) <= inputs(264) xor inputs(266) xor inputs(268) xor inputs(270) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(638) <= inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(639) <= inputs(505) xor inputs(507) xor inputs(509) xor inputs(511) ;
outputs(640) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(271) xor inputs(273) xor inputs(275) xor inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(641) <= inputs(127) xor inputs(129) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(271) xor inputs(273) xor inputs(275) xor inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(642) <= inputs(15) xor inputs(17) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(271) xor inputs(273) xor inputs(275) xor inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(643) <= inputs(271) xor inputs(273) xor inputs(275) xor inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(644) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(166) xor inputs(168) xor inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(645) <= inputs(166) xor inputs(168) xor inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(646) <= inputs(38) xor inputs(39) xor inputs(42) xor inputs(44) xor inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(647) <= inputs(389) xor inputs(391) xor inputs(397) xor inputs(399) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(648) <= inputs(1) xor inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(17) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(649) <= inputs(132) xor inputs(133) xor inputs(138) xor inputs(140) xor inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(650) <= inputs(17) xor inputs(19) xor inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(651) <= inputs(325) xor inputs(327) xor inputs(333) xor inputs(335) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(652) <= inputs(1) xor inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(653) <= inputs(212) xor inputs(214) xor inputs(220) xor inputs(222) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(654) <= inputs(69) xor inputs(71) xor inputs(76) xor inputs(78) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(655) <= inputs(453) xor inputs(455) xor inputs(461) xor inputs(463) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(656) <= inputs(0) xor inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(131) xor inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(657) <= inputs(127) xor inputs(129) xor inputs(131) xor inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(658) <= inputs(15) xor inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(659) <= inputs(294) xor inputs(296) xor inputs(302) xor inputs(304) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(660) <= inputs(0) xor inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(661) <= inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(662) <= inputs(45) xor inputs(50) xor inputs(52) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(663) <= inputs(421) xor inputs(423) xor inputs(429) xor inputs(431) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(664) <= inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(665) <= inputs(141) xor inputs(143) xor inputs(148) xor inputs(150) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(666) <= inputs(20) xor inputs(22) xor inputs(24) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(667) <= inputs(357) xor inputs(359) xor inputs(365) xor inputs(367) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(668) <= inputs(3) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(669) <= inputs(244) xor inputs(246) xor inputs(252) xor inputs(254) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(670) <= inputs(100) xor inputs(102) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(671) <= inputs(485) xor inputs(487) xor inputs(493) xor inputs(495) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(672) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(19) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(39) xor inputs(42) xor inputs(44) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(131) xor inputs(133) xor inputs(138) xor inputs(140) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(673) <= inputs(127) xor inputs(129) xor inputs(131) xor inputs(133) xor inputs(138) xor inputs(140) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(674) <= inputs(15) xor inputs(17) xor inputs(19) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(39) xor inputs(42) xor inputs(44) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(675) <= inputs(279) xor inputs(281) xor inputs(287) xor inputs(289) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(676) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(39) xor inputs(42) xor inputs(44) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(677) <= inputs(170) xor inputs(172) xor inputs(177) xor inputs(179) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(678) <= inputs(39) xor inputs(42) xor inputs(44) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(679) <= inputs(405) xor inputs(407) xor inputs(413) xor inputs(415) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(680) <= inputs(1) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(17) xor inputs(19) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(133) xor inputs(138) xor inputs(140) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(681) <= inputs(133) xor inputs(138) xor inputs(140) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(682) <= inputs(17) xor inputs(19) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(683) <= inputs(341) xor inputs(343) xor inputs(349) xor inputs(351) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(684) <= inputs(1) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(685) <= inputs(228) xor inputs(230) xor inputs(236) xor inputs(238) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(686) <= inputs(84) xor inputs(86) xor inputs(92) xor inputs(94) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(687) <= inputs(469) xor inputs(471) xor inputs(477) xor inputs(479) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(688) <= inputs(0) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(127) xor inputs(129) xor inputs(131) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(689) <= inputs(127) xor inputs(129) xor inputs(131) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(690) <= inputs(15) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(691) <= inputs(310) xor inputs(312) xor inputs(318) xor inputs(320) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(692) <= inputs(0) xor inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(693) <= inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(694) <= inputs(57) xor inputs(59) xor inputs(65) xor inputs(67) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(695) <= inputs(437) xor inputs(439) xor inputs(445) xor inputs(447) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(696) <= inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(697) <= inputs(155) xor inputs(157) xor inputs(163) xor inputs(165) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(698) <= inputs(27) xor inputs(29) xor inputs(35) xor inputs(37) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(699) <= inputs(373) xor inputs(375) xor inputs(381) xor inputs(383) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(700) <= inputs(5) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(701) <= inputs(260) xor inputs(262) xor inputs(268) xor inputs(270) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(702) <= inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(703) <= inputs(501) xor inputs(503) xor inputs(509) xor inputs(511) ;
outputs(704) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(19) xor inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(42) xor inputs(44) xor inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(129) xor inputs(131) xor inputs(132) xor inputs(138) xor inputs(140) xor inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(177) xor inputs(179) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(273) xor inputs(275) xor inputs(287) xor inputs(289) xor inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(705) <= inputs(129) xor inputs(131) xor inputs(132) xor inputs(138) xor inputs(140) xor inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(166) xor inputs(168) xor inputs(177) xor inputs(179) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(273) xor inputs(275) xor inputs(287) xor inputs(289) xor inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(706) <= inputs(15) xor inputs(17) xor inputs(19) xor inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(38) xor inputs(42) xor inputs(44) xor inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(273) xor inputs(275) xor inputs(287) xor inputs(289) xor inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(707) <= inputs(273) xor inputs(275) xor inputs(287) xor inputs(289) xor inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(708) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(12) xor inputs(14) xor inputs(38) xor inputs(42) xor inputs(44) xor inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(166) xor inputs(168) xor inputs(177) xor inputs(179) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(709) <= inputs(166) xor inputs(168) xor inputs(177) xor inputs(179) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(710) <= inputs(38) xor inputs(42) xor inputs(44) xor inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(711) <= inputs(397) xor inputs(399) xor inputs(413) xor inputs(415) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(712) <= inputs(1) xor inputs(3) xor inputs(12) xor inputs(14) xor inputs(17) xor inputs(19) xor inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(138) xor inputs(140) xor inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(713) <= inputs(132) xor inputs(138) xor inputs(140) xor inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(714) <= inputs(17) xor inputs(19) xor inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(715) <= inputs(333) xor inputs(335) xor inputs(349) xor inputs(351) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(716) <= inputs(1) xor inputs(3) xor inputs(12) xor inputs(14) xor inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(717) <= inputs(220) xor inputs(222) xor inputs(236) xor inputs(238) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(718) <= inputs(76) xor inputs(78) xor inputs(92) xor inputs(94) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(719) <= inputs(461) xor inputs(463) xor inputs(477) xor inputs(479) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(720) <= inputs(0) xor inputs(3) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(129) xor inputs(131) xor inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(721) <= inputs(129) xor inputs(131) xor inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(722) <= inputs(15) xor inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(723) <= inputs(302) xor inputs(304) xor inputs(318) xor inputs(320) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(724) <= inputs(0) xor inputs(3) xor inputs(12) xor inputs(14) xor inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(725) <= inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(726) <= inputs(50) xor inputs(52) xor inputs(65) xor inputs(67) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(727) <= inputs(429) xor inputs(431) xor inputs(445) xor inputs(447) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(728) <= inputs(3) xor inputs(12) xor inputs(14) xor inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(729) <= inputs(148) xor inputs(150) xor inputs(163) xor inputs(165) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(730) <= inputs(22) xor inputs(24) xor inputs(35) xor inputs(37) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(731) <= inputs(365) xor inputs(367) xor inputs(381) xor inputs(383) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(732) <= inputs(3) xor inputs(12) xor inputs(14) xor inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(733) <= inputs(252) xor inputs(254) xor inputs(268) xor inputs(270) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(734) <= inputs(108) xor inputs(110) xor inputs(124) xor inputs(126) xor inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(735) <= inputs(493) xor inputs(495) xor inputs(509) xor inputs(511) ;
outputs(736) <= inputs(0) xor inputs(1) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(17) xor inputs(19) xor inputs(35) xor inputs(37) xor inputs(42) xor inputs(44) xor inputs(65) xor inputs(67) xor inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(129) xor inputs(131) xor inputs(138) xor inputs(140) xor inputs(163) xor inputs(165) xor inputs(177) xor inputs(179) xor inputs(205) xor inputs(207) xor inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(287) xor inputs(289) xor inputs(318) xor inputs(320) xor inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(737) <= inputs(129) xor inputs(131) xor inputs(138) xor inputs(140) xor inputs(163) xor inputs(165) xor inputs(177) xor inputs(179) xor inputs(205) xor inputs(207) xor inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(287) xor inputs(289) xor inputs(318) xor inputs(320) xor inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(738) <= inputs(15) xor inputs(17) xor inputs(19) xor inputs(35) xor inputs(37) xor inputs(42) xor inputs(44) xor inputs(65) xor inputs(67) xor inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(287) xor inputs(289) xor inputs(318) xor inputs(320) xor inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(739) <= inputs(287) xor inputs(289) xor inputs(318) xor inputs(320) xor inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(740) <= inputs(0) xor inputs(1) xor inputs(12) xor inputs(14) xor inputs(42) xor inputs(44) xor inputs(65) xor inputs(67) xor inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(177) xor inputs(179) xor inputs(205) xor inputs(207) xor inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(741) <= inputs(177) xor inputs(179) xor inputs(205) xor inputs(207) xor inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(742) <= inputs(42) xor inputs(44) xor inputs(65) xor inputs(67) xor inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(743) <= inputs(413) xor inputs(415) xor inputs(445) xor inputs(447) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(744) <= inputs(1) xor inputs(12) xor inputs(14) xor inputs(17) xor inputs(19) xor inputs(35) xor inputs(37) xor inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(138) xor inputs(140) xor inputs(163) xor inputs(165) xor inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(745) <= inputs(138) xor inputs(140) xor inputs(163) xor inputs(165) xor inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(746) <= inputs(17) xor inputs(19) xor inputs(35) xor inputs(37) xor inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(747) <= inputs(349) xor inputs(351) xor inputs(381) xor inputs(383) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(748) <= inputs(1) xor inputs(12) xor inputs(14) xor inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(749) <= inputs(236) xor inputs(238) xor inputs(268) xor inputs(270) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(750) <= inputs(92) xor inputs(94) xor inputs(124) xor inputs(126) xor inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(751) <= inputs(477) xor inputs(479) xor inputs(509) xor inputs(511) ;
outputs(752) <= inputs(0) xor inputs(12) xor inputs(14) xor inputs(15) xor inputs(35) xor inputs(37) xor inputs(65) xor inputs(67) xor inputs(124) xor inputs(126) xor inputs(129) xor inputs(131) xor inputs(163) xor inputs(165) xor inputs(205) xor inputs(207) xor inputs(268) xor inputs(270) xor inputs(318) xor inputs(320) xor inputs(381) xor inputs(383) xor inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(753) <= inputs(129) xor inputs(131) xor inputs(163) xor inputs(165) xor inputs(205) xor inputs(207) xor inputs(268) xor inputs(270) xor inputs(318) xor inputs(320) xor inputs(381) xor inputs(383) xor inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(754) <= inputs(15) xor inputs(35) xor inputs(37) xor inputs(65) xor inputs(67) xor inputs(124) xor inputs(126) xor inputs(318) xor inputs(320) xor inputs(381) xor inputs(383) xor inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(755) <= inputs(318) xor inputs(320) xor inputs(381) xor inputs(383) xor inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(756) <= inputs(0) xor inputs(12) xor inputs(14) xor inputs(65) xor inputs(67) xor inputs(124) xor inputs(126) xor inputs(205) xor inputs(207) xor inputs(268) xor inputs(270) xor inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(757) <= inputs(205) xor inputs(207) xor inputs(268) xor inputs(270) xor inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(758) <= inputs(65) xor inputs(67) xor inputs(124) xor inputs(126) xor inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(759) <= inputs(445) xor inputs(447) xor inputs(509) xor inputs(511) ;
outputs(760) <= inputs(12) xor inputs(14) xor inputs(35) xor inputs(37) xor inputs(124) xor inputs(126) xor inputs(163) xor inputs(165) xor inputs(268) xor inputs(270) xor inputs(381) xor inputs(383) xor inputs(509) xor inputs(511) ;
outputs(761) <= inputs(163) xor inputs(165) xor inputs(268) xor inputs(270) xor inputs(381) xor inputs(383) xor inputs(509) xor inputs(511) ;
outputs(762) <= inputs(35) xor inputs(37) xor inputs(124) xor inputs(126) xor inputs(381) xor inputs(383) xor inputs(509) xor inputs(511) ;
outputs(763) <= inputs(381) xor inputs(383) xor inputs(509) xor inputs(511) ;
outputs(764) <= inputs(12) xor inputs(14) xor inputs(124) xor inputs(126) xor inputs(268) xor inputs(270) xor inputs(509) xor inputs(511) ;
outputs(765) <= inputs(268) xor inputs(270) xor inputs(509) xor inputs(511) ;
outputs(766) <= inputs(124) xor inputs(126) xor inputs(509) xor inputs(511) ;
outputs(767) <= inputs(509) xor inputs(511) ;
outputs(768) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(44) xor inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(136) xor inputs(140) xor inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(168) xor inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(275) xor inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(769) <= inputs(127) xor inputs(128) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(136) xor inputs(140) xor inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(168) xor inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(271) xor inputs(272) xor inputs(275) xor inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(770) <= inputs(15) xor inputs(16) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(44) xor inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(271) xor inputs(272) xor inputs(275) xor inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(771) <= inputs(271) xor inputs(272) xor inputs(275) xor inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(772) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(44) xor inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(168) xor inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(773) <= inputs(168) xor inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(774) <= inputs(38) xor inputs(39) xor inputs(40) xor inputs(44) xor inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(775) <= inputs(387) xor inputs(391) xor inputs(395) xor inputs(399) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(776) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(16) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(136) xor inputs(140) xor inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(777) <= inputs(132) xor inputs(133) xor inputs(136) xor inputs(140) xor inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(778) <= inputs(16) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(779) <= inputs(323) xor inputs(327) xor inputs(331) xor inputs(335) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(780) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(781) <= inputs(210) xor inputs(214) xor inputs(218) xor inputs(222) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(782) <= inputs(68) xor inputs(71) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(783) <= inputs(451) xor inputs(455) xor inputs(459) xor inputs(463) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(784) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(131) xor inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(785) <= inputs(127) xor inputs(128) xor inputs(131) xor inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(786) <= inputs(15) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(787) <= inputs(292) xor inputs(296) xor inputs(300) xor inputs(304) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(788) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(789) <= inputs(180) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(790) <= inputs(45) xor inputs(48) xor inputs(52) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(791) <= inputs(419) xor inputs(423) xor inputs(427) xor inputs(431) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(792) <= inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(793) <= inputs(143) xor inputs(146) xor inputs(150) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(794) <= inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(795) <= inputs(355) xor inputs(359) xor inputs(363) xor inputs(367) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(796) <= inputs(3) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(797) <= inputs(242) xor inputs(246) xor inputs(250) xor inputs(254) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(798) <= inputs(98) xor inputs(102) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(799) <= inputs(483) xor inputs(487) xor inputs(491) xor inputs(495) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(800) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(19) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(44) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(131) xor inputs(133) xor inputs(136) xor inputs(140) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(801) <= inputs(127) xor inputs(128) xor inputs(131) xor inputs(133) xor inputs(136) xor inputs(140) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(802) <= inputs(15) xor inputs(16) xor inputs(19) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(39) xor inputs(40) xor inputs(44) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(803) <= inputs(277) xor inputs(281) xor inputs(285) xor inputs(289) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(804) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(39) xor inputs(40) xor inputs(44) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(805) <= inputs(169) xor inputs(172) xor inputs(175) xor inputs(179) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(806) <= inputs(39) xor inputs(40) xor inputs(44) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(807) <= inputs(403) xor inputs(407) xor inputs(411) xor inputs(415) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(808) <= inputs(1) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(16) xor inputs(19) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(133) xor inputs(136) xor inputs(140) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(809) <= inputs(133) xor inputs(136) xor inputs(140) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(810) <= inputs(16) xor inputs(19) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(811) <= inputs(339) xor inputs(343) xor inputs(347) xor inputs(351) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(812) <= inputs(1) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(813) <= inputs(226) xor inputs(230) xor inputs(234) xor inputs(238) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(814) <= inputs(82) xor inputs(86) xor inputs(90) xor inputs(94) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(815) <= inputs(467) xor inputs(471) xor inputs(475) xor inputs(479) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(816) <= inputs(0) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(131) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(817) <= inputs(127) xor inputs(128) xor inputs(131) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(818) <= inputs(15) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(819) <= inputs(308) xor inputs(312) xor inputs(316) xor inputs(320) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(820) <= inputs(0) xor inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(821) <= inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(822) <= inputs(55) xor inputs(59) xor inputs(63) xor inputs(67) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(823) <= inputs(435) xor inputs(439) xor inputs(443) xor inputs(447) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(824) <= inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(825) <= inputs(153) xor inputs(157) xor inputs(161) xor inputs(165) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(826) <= inputs(25) xor inputs(29) xor inputs(33) xor inputs(37) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(827) <= inputs(371) xor inputs(375) xor inputs(379) xor inputs(383) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(828) <= inputs(4) xor inputs(7) xor inputs(10) xor inputs(14) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(829) <= inputs(258) xor inputs(262) xor inputs(266) xor inputs(270) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(830) <= inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(831) <= inputs(499) xor inputs(503) xor inputs(507) xor inputs(511) ;
outputs(832) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(19) xor inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(44) xor inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(128) xor inputs(131) xor inputs(132) xor inputs(136) xor inputs(140) xor inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(168) xor inputs(175) xor inputs(179) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(272) xor inputs(275) xor inputs(285) xor inputs(289) xor inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(833) <= inputs(128) xor inputs(131) xor inputs(132) xor inputs(136) xor inputs(140) xor inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(168) xor inputs(175) xor inputs(179) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(272) xor inputs(275) xor inputs(285) xor inputs(289) xor inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(834) <= inputs(15) xor inputs(16) xor inputs(19) xor inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(40) xor inputs(44) xor inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(272) xor inputs(275) xor inputs(285) xor inputs(289) xor inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(835) <= inputs(272) xor inputs(275) xor inputs(285) xor inputs(289) xor inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(836) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(10) xor inputs(14) xor inputs(38) xor inputs(40) xor inputs(44) xor inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(168) xor inputs(175) xor inputs(179) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(837) <= inputs(168) xor inputs(175) xor inputs(179) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(838) <= inputs(38) xor inputs(40) xor inputs(44) xor inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(839) <= inputs(395) xor inputs(399) xor inputs(411) xor inputs(415) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(840) <= inputs(1) xor inputs(3) xor inputs(10) xor inputs(14) xor inputs(16) xor inputs(19) xor inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(132) xor inputs(136) xor inputs(140) xor inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(841) <= inputs(132) xor inputs(136) xor inputs(140) xor inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(842) <= inputs(16) xor inputs(19) xor inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(843) <= inputs(331) xor inputs(335) xor inputs(347) xor inputs(351) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(844) <= inputs(1) xor inputs(3) xor inputs(10) xor inputs(14) xor inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(845) <= inputs(218) xor inputs(222) xor inputs(234) xor inputs(238) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(846) <= inputs(74) xor inputs(78) xor inputs(90) xor inputs(94) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(847) <= inputs(459) xor inputs(463) xor inputs(475) xor inputs(479) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(848) <= inputs(0) xor inputs(3) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(128) xor inputs(131) xor inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(849) <= inputs(128) xor inputs(131) xor inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(850) <= inputs(15) xor inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(851) <= inputs(300) xor inputs(304) xor inputs(316) xor inputs(320) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(852) <= inputs(0) xor inputs(3) xor inputs(10) xor inputs(14) xor inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(853) <= inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(854) <= inputs(48) xor inputs(52) xor inputs(63) xor inputs(67) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(855) <= inputs(427) xor inputs(431) xor inputs(443) xor inputs(447) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(856) <= inputs(3) xor inputs(10) xor inputs(14) xor inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(857) <= inputs(146) xor inputs(150) xor inputs(161) xor inputs(165) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(858) <= inputs(21) xor inputs(24) xor inputs(33) xor inputs(37) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(859) <= inputs(363) xor inputs(367) xor inputs(379) xor inputs(383) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(860) <= inputs(3) xor inputs(10) xor inputs(14) xor inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(861) <= inputs(250) xor inputs(254) xor inputs(266) xor inputs(270) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(862) <= inputs(106) xor inputs(110) xor inputs(122) xor inputs(126) xor inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(863) <= inputs(491) xor inputs(495) xor inputs(507) xor inputs(511) ;
outputs(864) <= inputs(0) xor inputs(1) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(19) xor inputs(33) xor inputs(37) xor inputs(40) xor inputs(44) xor inputs(63) xor inputs(67) xor inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(128) xor inputs(131) xor inputs(136) xor inputs(140) xor inputs(161) xor inputs(165) xor inputs(175) xor inputs(179) xor inputs(203) xor inputs(207) xor inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(285) xor inputs(289) xor inputs(316) xor inputs(320) xor inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(865) <= inputs(128) xor inputs(131) xor inputs(136) xor inputs(140) xor inputs(161) xor inputs(165) xor inputs(175) xor inputs(179) xor inputs(203) xor inputs(207) xor inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(285) xor inputs(289) xor inputs(316) xor inputs(320) xor inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(866) <= inputs(15) xor inputs(16) xor inputs(19) xor inputs(33) xor inputs(37) xor inputs(40) xor inputs(44) xor inputs(63) xor inputs(67) xor inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(285) xor inputs(289) xor inputs(316) xor inputs(320) xor inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(867) <= inputs(285) xor inputs(289) xor inputs(316) xor inputs(320) xor inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(868) <= inputs(0) xor inputs(1) xor inputs(10) xor inputs(14) xor inputs(40) xor inputs(44) xor inputs(63) xor inputs(67) xor inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(175) xor inputs(179) xor inputs(203) xor inputs(207) xor inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(869) <= inputs(175) xor inputs(179) xor inputs(203) xor inputs(207) xor inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(870) <= inputs(40) xor inputs(44) xor inputs(63) xor inputs(67) xor inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(871) <= inputs(411) xor inputs(415) xor inputs(443) xor inputs(447) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(872) <= inputs(1) xor inputs(10) xor inputs(14) xor inputs(16) xor inputs(19) xor inputs(33) xor inputs(37) xor inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(136) xor inputs(140) xor inputs(161) xor inputs(165) xor inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(873) <= inputs(136) xor inputs(140) xor inputs(161) xor inputs(165) xor inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(874) <= inputs(16) xor inputs(19) xor inputs(33) xor inputs(37) xor inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(875) <= inputs(347) xor inputs(351) xor inputs(379) xor inputs(383) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(876) <= inputs(1) xor inputs(10) xor inputs(14) xor inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(877) <= inputs(234) xor inputs(238) xor inputs(266) xor inputs(270) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(878) <= inputs(90) xor inputs(94) xor inputs(122) xor inputs(126) xor inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(879) <= inputs(475) xor inputs(479) xor inputs(507) xor inputs(511) ;
outputs(880) <= inputs(0) xor inputs(10) xor inputs(14) xor inputs(15) xor inputs(33) xor inputs(37) xor inputs(63) xor inputs(67) xor inputs(122) xor inputs(126) xor inputs(128) xor inputs(131) xor inputs(161) xor inputs(165) xor inputs(203) xor inputs(207) xor inputs(266) xor inputs(270) xor inputs(316) xor inputs(320) xor inputs(379) xor inputs(383) xor inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(881) <= inputs(128) xor inputs(131) xor inputs(161) xor inputs(165) xor inputs(203) xor inputs(207) xor inputs(266) xor inputs(270) xor inputs(316) xor inputs(320) xor inputs(379) xor inputs(383) xor inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(882) <= inputs(15) xor inputs(33) xor inputs(37) xor inputs(63) xor inputs(67) xor inputs(122) xor inputs(126) xor inputs(316) xor inputs(320) xor inputs(379) xor inputs(383) xor inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(883) <= inputs(316) xor inputs(320) xor inputs(379) xor inputs(383) xor inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(884) <= inputs(0) xor inputs(10) xor inputs(14) xor inputs(63) xor inputs(67) xor inputs(122) xor inputs(126) xor inputs(203) xor inputs(207) xor inputs(266) xor inputs(270) xor inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(885) <= inputs(203) xor inputs(207) xor inputs(266) xor inputs(270) xor inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(886) <= inputs(63) xor inputs(67) xor inputs(122) xor inputs(126) xor inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(887) <= inputs(443) xor inputs(447) xor inputs(507) xor inputs(511) ;
outputs(888) <= inputs(10) xor inputs(14) xor inputs(33) xor inputs(37) xor inputs(122) xor inputs(126) xor inputs(161) xor inputs(165) xor inputs(266) xor inputs(270) xor inputs(379) xor inputs(383) xor inputs(507) xor inputs(511) ;
outputs(889) <= inputs(161) xor inputs(165) xor inputs(266) xor inputs(270) xor inputs(379) xor inputs(383) xor inputs(507) xor inputs(511) ;
outputs(890) <= inputs(33) xor inputs(37) xor inputs(122) xor inputs(126) xor inputs(379) xor inputs(383) xor inputs(507) xor inputs(511) ;
outputs(891) <= inputs(379) xor inputs(383) xor inputs(507) xor inputs(511) ;
outputs(892) <= inputs(10) xor inputs(14) xor inputs(122) xor inputs(126) xor inputs(266) xor inputs(270) xor inputs(507) xor inputs(511) ;
outputs(893) <= inputs(266) xor inputs(270) xor inputs(507) xor inputs(511) ;
outputs(894) <= inputs(122) xor inputs(126) xor inputs(507) xor inputs(511) ;
outputs(895) <= inputs(507) xor inputs(511) ;
outputs(896) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(7) xor inputs(14) xor inputs(15) xor inputs(19) xor inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(44) xor inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(127) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(140) xor inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(168) xor inputs(172) xor inputs(179) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(271) xor inputs(275) xor inputs(281) xor inputs(289) xor inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(897) <= inputs(127) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(140) xor inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(168) xor inputs(172) xor inputs(179) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(271) xor inputs(275) xor inputs(281) xor inputs(289) xor inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(898) <= inputs(15) xor inputs(19) xor inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(44) xor inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(271) xor inputs(275) xor inputs(281) xor inputs(289) xor inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(899) <= inputs(271) xor inputs(275) xor inputs(281) xor inputs(289) xor inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(900) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(7) xor inputs(14) xor inputs(38) xor inputs(39) xor inputs(44) xor inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(168) xor inputs(172) xor inputs(179) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(901) <= inputs(168) xor inputs(172) xor inputs(179) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(902) <= inputs(38) xor inputs(39) xor inputs(44) xor inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(903) <= inputs(391) xor inputs(399) xor inputs(407) xor inputs(415) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(904) <= inputs(1) xor inputs(3) xor inputs(7) xor inputs(14) xor inputs(19) xor inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(132) xor inputs(133) xor inputs(140) xor inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(905) <= inputs(132) xor inputs(133) xor inputs(140) xor inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(906) <= inputs(19) xor inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(907) <= inputs(327) xor inputs(335) xor inputs(343) xor inputs(351) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(908) <= inputs(1) xor inputs(3) xor inputs(7) xor inputs(14) xor inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(909) <= inputs(214) xor inputs(222) xor inputs(230) xor inputs(238) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(910) <= inputs(71) xor inputs(78) xor inputs(86) xor inputs(94) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(911) <= inputs(455) xor inputs(463) xor inputs(471) xor inputs(479) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(912) <= inputs(0) xor inputs(3) xor inputs(7) xor inputs(14) xor inputs(15) xor inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(127) xor inputs(131) xor inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(913) <= inputs(127) xor inputs(131) xor inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(914) <= inputs(15) xor inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(915) <= inputs(296) xor inputs(304) xor inputs(312) xor inputs(320) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(916) <= inputs(0) xor inputs(3) xor inputs(7) xor inputs(14) xor inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(917) <= inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(918) <= inputs(45) xor inputs(52) xor inputs(59) xor inputs(67) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(919) <= inputs(423) xor inputs(431) xor inputs(439) xor inputs(447) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(920) <= inputs(3) xor inputs(7) xor inputs(14) xor inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(921) <= inputs(143) xor inputs(150) xor inputs(157) xor inputs(165) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(922) <= inputs(20) xor inputs(24) xor inputs(29) xor inputs(37) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(923) <= inputs(359) xor inputs(367) xor inputs(375) xor inputs(383) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(924) <= inputs(3) xor inputs(7) xor inputs(14) xor inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(925) <= inputs(246) xor inputs(254) xor inputs(262) xor inputs(270) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(926) <= inputs(102) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(927) <= inputs(487) xor inputs(495) xor inputs(503) xor inputs(511) ;
outputs(928) <= inputs(0) xor inputs(1) xor inputs(7) xor inputs(14) xor inputs(15) xor inputs(19) xor inputs(29) xor inputs(37) xor inputs(39) xor inputs(44) xor inputs(59) xor inputs(67) xor inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(127) xor inputs(131) xor inputs(133) xor inputs(140) xor inputs(157) xor inputs(165) xor inputs(172) xor inputs(179) xor inputs(199) xor inputs(207) xor inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(281) xor inputs(289) xor inputs(312) xor inputs(320) xor inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(929) <= inputs(127) xor inputs(131) xor inputs(133) xor inputs(140) xor inputs(157) xor inputs(165) xor inputs(172) xor inputs(179) xor inputs(199) xor inputs(207) xor inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(281) xor inputs(289) xor inputs(312) xor inputs(320) xor inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(930) <= inputs(15) xor inputs(19) xor inputs(29) xor inputs(37) xor inputs(39) xor inputs(44) xor inputs(59) xor inputs(67) xor inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(281) xor inputs(289) xor inputs(312) xor inputs(320) xor inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(931) <= inputs(281) xor inputs(289) xor inputs(312) xor inputs(320) xor inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(932) <= inputs(0) xor inputs(1) xor inputs(7) xor inputs(14) xor inputs(39) xor inputs(44) xor inputs(59) xor inputs(67) xor inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(172) xor inputs(179) xor inputs(199) xor inputs(207) xor inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(933) <= inputs(172) xor inputs(179) xor inputs(199) xor inputs(207) xor inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(934) <= inputs(39) xor inputs(44) xor inputs(59) xor inputs(67) xor inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(935) <= inputs(407) xor inputs(415) xor inputs(439) xor inputs(447) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(936) <= inputs(1) xor inputs(7) xor inputs(14) xor inputs(19) xor inputs(29) xor inputs(37) xor inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(133) xor inputs(140) xor inputs(157) xor inputs(165) xor inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(937) <= inputs(133) xor inputs(140) xor inputs(157) xor inputs(165) xor inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(938) <= inputs(19) xor inputs(29) xor inputs(37) xor inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(939) <= inputs(343) xor inputs(351) xor inputs(375) xor inputs(383) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(940) <= inputs(1) xor inputs(7) xor inputs(14) xor inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(941) <= inputs(230) xor inputs(238) xor inputs(262) xor inputs(270) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(942) <= inputs(86) xor inputs(94) xor inputs(118) xor inputs(126) xor inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(943) <= inputs(471) xor inputs(479) xor inputs(503) xor inputs(511) ;
outputs(944) <= inputs(0) xor inputs(7) xor inputs(14) xor inputs(15) xor inputs(29) xor inputs(37) xor inputs(59) xor inputs(67) xor inputs(118) xor inputs(126) xor inputs(127) xor inputs(131) xor inputs(157) xor inputs(165) xor inputs(199) xor inputs(207) xor inputs(262) xor inputs(270) xor inputs(312) xor inputs(320) xor inputs(375) xor inputs(383) xor inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(945) <= inputs(127) xor inputs(131) xor inputs(157) xor inputs(165) xor inputs(199) xor inputs(207) xor inputs(262) xor inputs(270) xor inputs(312) xor inputs(320) xor inputs(375) xor inputs(383) xor inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(946) <= inputs(15) xor inputs(29) xor inputs(37) xor inputs(59) xor inputs(67) xor inputs(118) xor inputs(126) xor inputs(312) xor inputs(320) xor inputs(375) xor inputs(383) xor inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(947) <= inputs(312) xor inputs(320) xor inputs(375) xor inputs(383) xor inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(948) <= inputs(0) xor inputs(7) xor inputs(14) xor inputs(59) xor inputs(67) xor inputs(118) xor inputs(126) xor inputs(199) xor inputs(207) xor inputs(262) xor inputs(270) xor inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(949) <= inputs(199) xor inputs(207) xor inputs(262) xor inputs(270) xor inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(950) <= inputs(59) xor inputs(67) xor inputs(118) xor inputs(126) xor inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(951) <= inputs(439) xor inputs(447) xor inputs(503) xor inputs(511) ;
outputs(952) <= inputs(7) xor inputs(14) xor inputs(29) xor inputs(37) xor inputs(118) xor inputs(126) xor inputs(157) xor inputs(165) xor inputs(262) xor inputs(270) xor inputs(375) xor inputs(383) xor inputs(503) xor inputs(511) ;
outputs(953) <= inputs(157) xor inputs(165) xor inputs(262) xor inputs(270) xor inputs(375) xor inputs(383) xor inputs(503) xor inputs(511) ;
outputs(954) <= inputs(29) xor inputs(37) xor inputs(118) xor inputs(126) xor inputs(375) xor inputs(383) xor inputs(503) xor inputs(511) ;
outputs(955) <= inputs(375) xor inputs(383) xor inputs(503) xor inputs(511) ;
outputs(956) <= inputs(7) xor inputs(14) xor inputs(118) xor inputs(126) xor inputs(262) xor inputs(270) xor inputs(503) xor inputs(511) ;
outputs(957) <= inputs(262) xor inputs(270) xor inputs(503) xor inputs(511) ;
outputs(958) <= inputs(118) xor inputs(126) xor inputs(503) xor inputs(511) ;
outputs(959) <= inputs(503) xor inputs(511) ;
outputs(960) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(14) xor inputs(15) xor inputs(19) xor inputs(24) xor inputs(37) xor inputs(38) xor inputs(44) xor inputs(52) xor inputs(67) xor inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(140) xor inputs(150) xor inputs(165) xor inputs(168) xor inputs(179) xor inputs(191) xor inputs(207) xor inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(275) xor inputs(289) xor inputs(304) xor inputs(320) xor inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(961) <= inputs(131) xor inputs(132) xor inputs(140) xor inputs(150) xor inputs(165) xor inputs(168) xor inputs(179) xor inputs(191) xor inputs(207) xor inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(275) xor inputs(289) xor inputs(304) xor inputs(320) xor inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(962) <= inputs(15) xor inputs(19) xor inputs(24) xor inputs(37) xor inputs(38) xor inputs(44) xor inputs(52) xor inputs(67) xor inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(275) xor inputs(289) xor inputs(304) xor inputs(320) xor inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(963) <= inputs(275) xor inputs(289) xor inputs(304) xor inputs(320) xor inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(964) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(14) xor inputs(38) xor inputs(44) xor inputs(52) xor inputs(67) xor inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(168) xor inputs(179) xor inputs(191) xor inputs(207) xor inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(965) <= inputs(168) xor inputs(179) xor inputs(191) xor inputs(207) xor inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(966) <= inputs(38) xor inputs(44) xor inputs(52) xor inputs(67) xor inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(967) <= inputs(399) xor inputs(415) xor inputs(431) xor inputs(447) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(968) <= inputs(1) xor inputs(3) xor inputs(14) xor inputs(19) xor inputs(24) xor inputs(37) xor inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(132) xor inputs(140) xor inputs(150) xor inputs(165) xor inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(969) <= inputs(132) xor inputs(140) xor inputs(150) xor inputs(165) xor inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(970) <= inputs(19) xor inputs(24) xor inputs(37) xor inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(971) <= inputs(335) xor inputs(351) xor inputs(367) xor inputs(383) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(972) <= inputs(1) xor inputs(3) xor inputs(14) xor inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(973) <= inputs(222) xor inputs(238) xor inputs(254) xor inputs(270) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(974) <= inputs(78) xor inputs(94) xor inputs(110) xor inputs(126) xor inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(975) <= inputs(463) xor inputs(479) xor inputs(495) xor inputs(511) ;
outputs(976) <= inputs(0) xor inputs(3) xor inputs(14) xor inputs(15) xor inputs(24) xor inputs(37) xor inputs(52) xor inputs(67) xor inputs(110) xor inputs(126) xor inputs(131) xor inputs(150) xor inputs(165) xor inputs(191) xor inputs(207) xor inputs(254) xor inputs(270) xor inputs(304) xor inputs(320) xor inputs(367) xor inputs(383) xor inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(977) <= inputs(131) xor inputs(150) xor inputs(165) xor inputs(191) xor inputs(207) xor inputs(254) xor inputs(270) xor inputs(304) xor inputs(320) xor inputs(367) xor inputs(383) xor inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(978) <= inputs(15) xor inputs(24) xor inputs(37) xor inputs(52) xor inputs(67) xor inputs(110) xor inputs(126) xor inputs(304) xor inputs(320) xor inputs(367) xor inputs(383) xor inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(979) <= inputs(304) xor inputs(320) xor inputs(367) xor inputs(383) xor inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(980) <= inputs(0) xor inputs(3) xor inputs(14) xor inputs(52) xor inputs(67) xor inputs(110) xor inputs(126) xor inputs(191) xor inputs(207) xor inputs(254) xor inputs(270) xor inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(981) <= inputs(191) xor inputs(207) xor inputs(254) xor inputs(270) xor inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(982) <= inputs(52) xor inputs(67) xor inputs(110) xor inputs(126) xor inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(983) <= inputs(431) xor inputs(447) xor inputs(495) xor inputs(511) ;
outputs(984) <= inputs(3) xor inputs(14) xor inputs(24) xor inputs(37) xor inputs(110) xor inputs(126) xor inputs(150) xor inputs(165) xor inputs(254) xor inputs(270) xor inputs(367) xor inputs(383) xor inputs(495) xor inputs(511) ;
outputs(985) <= inputs(150) xor inputs(165) xor inputs(254) xor inputs(270) xor inputs(367) xor inputs(383) xor inputs(495) xor inputs(511) ;
outputs(986) <= inputs(24) xor inputs(37) xor inputs(110) xor inputs(126) xor inputs(367) xor inputs(383) xor inputs(495) xor inputs(511) ;
outputs(987) <= inputs(367) xor inputs(383) xor inputs(495) xor inputs(511) ;
outputs(988) <= inputs(3) xor inputs(14) xor inputs(110) xor inputs(126) xor inputs(254) xor inputs(270) xor inputs(495) xor inputs(511) ;
outputs(989) <= inputs(254) xor inputs(270) xor inputs(495) xor inputs(511) ;
outputs(990) <= inputs(110) xor inputs(126) xor inputs(495) xor inputs(511) ;
outputs(991) <= inputs(495) xor inputs(511) ;
outputs(992) <= inputs(0) xor inputs(1) xor inputs(14) xor inputs(15) xor inputs(19) xor inputs(37) xor inputs(44) xor inputs(67) xor inputs(94) xor inputs(126) xor inputs(131) xor inputs(140) xor inputs(165) xor inputs(179) xor inputs(207) xor inputs(238) xor inputs(270) xor inputs(289) xor inputs(320) xor inputs(351) xor inputs(383) xor inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(993) <= inputs(131) xor inputs(140) xor inputs(165) xor inputs(179) xor inputs(207) xor inputs(238) xor inputs(270) xor inputs(289) xor inputs(320) xor inputs(351) xor inputs(383) xor inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(994) <= inputs(15) xor inputs(19) xor inputs(37) xor inputs(44) xor inputs(67) xor inputs(94) xor inputs(126) xor inputs(289) xor inputs(320) xor inputs(351) xor inputs(383) xor inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(995) <= inputs(289) xor inputs(320) xor inputs(351) xor inputs(383) xor inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(996) <= inputs(0) xor inputs(1) xor inputs(14) xor inputs(44) xor inputs(67) xor inputs(94) xor inputs(126) xor inputs(179) xor inputs(207) xor inputs(238) xor inputs(270) xor inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(997) <= inputs(179) xor inputs(207) xor inputs(238) xor inputs(270) xor inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(998) <= inputs(44) xor inputs(67) xor inputs(94) xor inputs(126) xor inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(999) <= inputs(415) xor inputs(447) xor inputs(479) xor inputs(511) ;
outputs(1000) <= inputs(1) xor inputs(14) xor inputs(19) xor inputs(37) xor inputs(94) xor inputs(126) xor inputs(140) xor inputs(165) xor inputs(238) xor inputs(270) xor inputs(351) xor inputs(383) xor inputs(479) xor inputs(511) ;
outputs(1001) <= inputs(140) xor inputs(165) xor inputs(238) xor inputs(270) xor inputs(351) xor inputs(383) xor inputs(479) xor inputs(511) ;
outputs(1002) <= inputs(19) xor inputs(37) xor inputs(94) xor inputs(126) xor inputs(351) xor inputs(383) xor inputs(479) xor inputs(511) ;
outputs(1003) <= inputs(351) xor inputs(383) xor inputs(479) xor inputs(511) ;
outputs(1004) <= inputs(1) xor inputs(14) xor inputs(94) xor inputs(126) xor inputs(238) xor inputs(270) xor inputs(479) xor inputs(511) ;
outputs(1005) <= inputs(238) xor inputs(270) xor inputs(479) xor inputs(511) ;
outputs(1006) <= inputs(94) xor inputs(126) xor inputs(479) xor inputs(511) ;
outputs(1007) <= inputs(479) xor inputs(511) ;
outputs(1008) <= inputs(0) xor inputs(14) xor inputs(15) xor inputs(37) xor inputs(67) xor inputs(126) xor inputs(131) xor inputs(165) xor inputs(207) xor inputs(270) xor inputs(320) xor inputs(383) xor inputs(447) xor inputs(511) ;
outputs(1009) <= inputs(131) xor inputs(165) xor inputs(207) xor inputs(270) xor inputs(320) xor inputs(383) xor inputs(447) xor inputs(511) ;
outputs(1010) <= inputs(15) xor inputs(37) xor inputs(67) xor inputs(126) xor inputs(320) xor inputs(383) xor inputs(447) xor inputs(511) ;
outputs(1011) <= inputs(320) xor inputs(383) xor inputs(447) xor inputs(511) ;
outputs(1012) <= inputs(0) xor inputs(14) xor inputs(67) xor inputs(126) xor inputs(207) xor inputs(270) xor inputs(447) xor inputs(511) ;
outputs(1013) <= inputs(207) xor inputs(270) xor inputs(447) xor inputs(511) ;
outputs(1014) <= inputs(67) xor inputs(126) xor inputs(447) xor inputs(511) ;
outputs(1015) <= inputs(447) xor inputs(511) ;
outputs(1016) <= inputs(14) xor inputs(37) xor inputs(126) xor inputs(165) xor inputs(270) xor inputs(383) xor inputs(511) ;
outputs(1017) <= inputs(165) xor inputs(270) xor inputs(383) xor inputs(511) ;
outputs(1018) <= inputs(37) xor inputs(126) xor inputs(383) xor inputs(511) ;
outputs(1019) <= inputs(383) xor inputs(511) ;
outputs(1020) <= inputs(14) xor inputs(126) xor inputs(270) xor inputs(511) ;
outputs(1021) <= inputs(270) xor inputs(511) ;
outputs(1022) <= inputs(126) xor inputs(511) ;
outputs(1023) <= inputs(511);

end Behavioral;


----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:13:37 04/03/2016 
-- Design Name: 
-- Module Name:    Encoder512 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.all;
use work.MyPackage.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Encoder512 is
	Port (inputs : in std_logic_vector(N/2-1 downto 0);
			outputs : out std_logic_vector(N-1 downto 0));
end Encoder512;

architecture Behavioral of Encoder512 is

begin

outputs(0) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(1) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(2) <= inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(3) <= inputs(135) xor inputs(136) xor inputs(137) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(4) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(5) <= inputs(83) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(6) <= inputs(19) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(7) <= inputs(192) xor inputs(193) xor inputs(194) xor inputs(195) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(8) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(9) <= inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(10) <= inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(11) <= inputs(160) xor inputs(161) xor inputs(162) xor inputs(163) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(12) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(13) <= inputs(104) xor inputs(105) xor inputs(106) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(14) <= inputs(34) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(15) <= inputs(224) xor inputs(225) xor inputs(226) xor inputs(227) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(16) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(17) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(18) <= inputs(7) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(19) <= inputs(145) xor inputs(146) xor inputs(147) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(20) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(21) <= inputs(89) xor inputs(90) xor inputs(91) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(22) <= inputs(22) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(23) <= inputs(208) xor inputs(209) xor inputs(210) xor inputs(211) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(24) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(25) <= inputs(70) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(26) <= inputs(9) xor inputs(10) xor inputs(11) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(27) <= inputs(176) xor inputs(177) xor inputs(178) xor inputs(179) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(28) <= inputs(1) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(29) <= inputs(119) xor inputs(120) xor inputs(121) xor inputs(122) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(30) <= inputs(47) xor inputs(48) xor inputs(49) xor inputs(50) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(31) <= inputs(240) xor inputs(241) xor inputs(242) xor inputs(243) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(32) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(33) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(34) <= inputs(7) xor inputs(8) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(35) <= inputs(138) xor inputs(139) xor inputs(140) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(36) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(37) <= inputs(84) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(38) <= inputs(19) xor inputs(20) xor inputs(21) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(39) <= inputs(200) xor inputs(201) xor inputs(202) xor inputs(203) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(40) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(41) <= inputs(66) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(42) <= inputs(8) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(43) <= inputs(168) xor inputs(169) xor inputs(170) xor inputs(171) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(44) <= inputs(0) xor inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(45) <= inputs(111) xor inputs(112) xor inputs(113) xor inputs(114) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(46) <= inputs(39) xor inputs(40) xor inputs(41) xor inputs(42) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(47) <= inputs(232) xor inputs(233) xor inputs(234) xor inputs(235) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(48) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(49) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(50) <= inputs(7) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(51) <= inputs(152) xor inputs(153) xor inputs(154) xor inputs(155) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(52) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(53) <= inputs(96) xor inputs(97) xor inputs(98) xor inputs(99) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(54) <= inputs(26) xor inputs(27) xor inputs(28) xor inputs(29) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(55) <= inputs(216) xor inputs(217) xor inputs(218) xor inputs(219) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(56) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(57) <= inputs(75) xor inputs(76) xor inputs(77) xor inputs(78) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(58) <= inputs(12) xor inputs(13) xor inputs(14) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(59) <= inputs(184) xor inputs(185) xor inputs(186) xor inputs(187) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(60) <= inputs(2) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(61) <= inputs(127) xor inputs(128) xor inputs(129) xor inputs(130) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(62) <= inputs(55) xor inputs(56) xor inputs(57) xor inputs(58) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(63) <= inputs(248) xor inputs(249) xor inputs(250) xor inputs(251) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(64) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(65) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(66) <= inputs(7) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(135) xor inputs(136) xor inputs(137) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(67) <= inputs(135) xor inputs(136) xor inputs(137) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(68) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(83) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(69) <= inputs(83) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(70) <= inputs(19) xor inputs(20) xor inputs(21) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(71) <= inputs(196) xor inputs(197) xor inputs(198) xor inputs(199) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(72) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(73) <= inputs(67) xor inputs(68) xor inputs(69) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(74) <= inputs(8) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(75) <= inputs(164) xor inputs(165) xor inputs(166) xor inputs(167) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(76) <= inputs(0) xor inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(77) <= inputs(107) xor inputs(108) xor inputs(109) xor inputs(110) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(78) <= inputs(35) xor inputs(36) xor inputs(37) xor inputs(38) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(79) <= inputs(228) xor inputs(229) xor inputs(230) xor inputs(231) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(80) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(81) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(82) <= inputs(7) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(83) <= inputs(148) xor inputs(149) xor inputs(150) xor inputs(151) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(84) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(85) <= inputs(92) xor inputs(93) xor inputs(94) xor inputs(95) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(86) <= inputs(23) xor inputs(24) xor inputs(25) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(87) <= inputs(212) xor inputs(213) xor inputs(214) xor inputs(215) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(88) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(89) <= inputs(71) xor inputs(72) xor inputs(73) xor inputs(74) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(90) <= inputs(9) xor inputs(10) xor inputs(11) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(91) <= inputs(180) xor inputs(181) xor inputs(182) xor inputs(183) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(92) <= inputs(1) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(93) <= inputs(123) xor inputs(124) xor inputs(125) xor inputs(126) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(94) <= inputs(51) xor inputs(52) xor inputs(53) xor inputs(54) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(95) <= inputs(244) xor inputs(245) xor inputs(246) xor inputs(247) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(96) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(97) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(98) <= inputs(7) xor inputs(8) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(99) <= inputs(141) xor inputs(142) xor inputs(143) xor inputs(144) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(100) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(19) xor inputs(20) xor inputs(21) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(101) <= inputs(85) xor inputs(86) xor inputs(87) xor inputs(88) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(102) <= inputs(19) xor inputs(20) xor inputs(21) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(103) <= inputs(204) xor inputs(205) xor inputs(206) xor inputs(207) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(104) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(67) xor inputs(68) xor inputs(69) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(105) <= inputs(67) xor inputs(68) xor inputs(69) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(106) <= inputs(8) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(107) <= inputs(172) xor inputs(173) xor inputs(174) xor inputs(175) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(108) <= inputs(0) xor inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(109) <= inputs(115) xor inputs(116) xor inputs(117) xor inputs(118) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(110) <= inputs(43) xor inputs(44) xor inputs(45) xor inputs(46) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(111) <= inputs(236) xor inputs(237) xor inputs(238) xor inputs(239) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(112) <= inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(63) xor inputs(64) xor inputs(65) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(113) <= inputs(63) xor inputs(64) xor inputs(65) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(114) <= inputs(7) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(115) <= inputs(156) xor inputs(157) xor inputs(158) xor inputs(159) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(116) <= inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(117) <= inputs(100) xor inputs(101) xor inputs(102) xor inputs(103) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(118) <= inputs(30) xor inputs(31) xor inputs(32) xor inputs(33) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(119) <= inputs(220) xor inputs(221) xor inputs(222) xor inputs(223) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(120) <= inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(121) <= inputs(79) xor inputs(80) xor inputs(81) xor inputs(82) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(122) <= inputs(15) xor inputs(16) xor inputs(17) xor inputs(18) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(123) <= inputs(188) xor inputs(189) xor inputs(190) xor inputs(191) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(124) <= inputs(3) xor inputs(4) xor inputs(5) xor inputs(6) xor inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(125) <= inputs(131) xor inputs(132) xor inputs(133) xor inputs(134) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(126) <= inputs(59) xor inputs(60) xor inputs(61) xor inputs(62) xor inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(127) <= inputs(252) xor inputs(253) xor inputs(254) xor inputs(255) ;
outputs(128) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(87) xor inputs(88) xor inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(137) xor inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(129) <= inputs(64) xor inputs(65) xor inputs(66) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(87) xor inputs(88) xor inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(137) xor inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(130) <= inputs(7) xor inputs(8) xor inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(136) xor inputs(137) xor inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(131) <= inputs(136) xor inputs(137) xor inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(132) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(83) xor inputs(84) xor inputs(87) xor inputs(88) xor inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(133) <= inputs(83) xor inputs(84) xor inputs(87) xor inputs(88) xor inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(134) <= inputs(20) xor inputs(21) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(135) <= inputs(194) xor inputs(195) xor inputs(198) xor inputs(199) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(136) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(66) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(137) <= inputs(66) xor inputs(68) xor inputs(69) xor inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(138) <= inputs(8) xor inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(139) <= inputs(162) xor inputs(163) xor inputs(166) xor inputs(167) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(140) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(141) <= inputs(105) xor inputs(106) xor inputs(109) xor inputs(110) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(142) <= inputs(34) xor inputs(37) xor inputs(38) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(143) <= inputs(226) xor inputs(227) xor inputs(230) xor inputs(231) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(144) <= inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(145) <= inputs(64) xor inputs(65) xor inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(146) <= inputs(7) xor inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(147) <= inputs(146) xor inputs(147) xor inputs(150) xor inputs(151) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(148) <= inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(149) <= inputs(90) xor inputs(91) xor inputs(94) xor inputs(95) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(150) <= inputs(22) xor inputs(24) xor inputs(25) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(151) <= inputs(210) xor inputs(211) xor inputs(214) xor inputs(215) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(152) <= inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(153) <= inputs(70) xor inputs(73) xor inputs(74) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(154) <= inputs(10) xor inputs(11) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(155) <= inputs(178) xor inputs(179) xor inputs(182) xor inputs(183) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(156) <= inputs(1) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(157) <= inputs(121) xor inputs(122) xor inputs(125) xor inputs(126) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(158) <= inputs(49) xor inputs(50) xor inputs(53) xor inputs(54) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(159) <= inputs(242) xor inputs(243) xor inputs(246) xor inputs(247) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(160) <= inputs(0) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(66) xor inputs(68) xor inputs(69) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(84) xor inputs(87) xor inputs(88) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(161) <= inputs(64) xor inputs(65) xor inputs(66) xor inputs(68) xor inputs(69) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(84) xor inputs(87) xor inputs(88) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(162) <= inputs(7) xor inputs(8) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(163) <= inputs(139) xor inputs(140) xor inputs(143) xor inputs(144) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(164) <= inputs(0) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(20) xor inputs(21) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(84) xor inputs(87) xor inputs(88) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(165) <= inputs(84) xor inputs(87) xor inputs(88) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(166) <= inputs(20) xor inputs(21) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(167) <= inputs(202) xor inputs(203) xor inputs(206) xor inputs(207) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(168) <= inputs(0) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(66) xor inputs(68) xor inputs(69) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(169) <= inputs(66) xor inputs(68) xor inputs(69) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(170) <= inputs(8) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(171) <= inputs(170) xor inputs(171) xor inputs(174) xor inputs(175) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(172) <= inputs(0) xor inputs(2) xor inputs(5) xor inputs(6) xor inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(173) <= inputs(113) xor inputs(114) xor inputs(117) xor inputs(118) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(174) <= inputs(41) xor inputs(42) xor inputs(45) xor inputs(46) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(175) <= inputs(234) xor inputs(235) xor inputs(238) xor inputs(239) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(176) <= inputs(2) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(177) <= inputs(64) xor inputs(65) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(178) <= inputs(7) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(179) <= inputs(154) xor inputs(155) xor inputs(158) xor inputs(159) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(180) <= inputs(2) xor inputs(5) xor inputs(6) xor inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(181) <= inputs(98) xor inputs(99) xor inputs(102) xor inputs(103) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(182) <= inputs(28) xor inputs(29) xor inputs(32) xor inputs(33) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(183) <= inputs(218) xor inputs(219) xor inputs(222) xor inputs(223) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(184) <= inputs(2) xor inputs(5) xor inputs(6) xor inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(185) <= inputs(77) xor inputs(78) xor inputs(81) xor inputs(82) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(186) <= inputs(13) xor inputs(14) xor inputs(17) xor inputs(18) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(187) <= inputs(186) xor inputs(187) xor inputs(190) xor inputs(191) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(188) <= inputs(2) xor inputs(5) xor inputs(6) xor inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(189) <= inputs(129) xor inputs(130) xor inputs(133) xor inputs(134) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(190) <= inputs(57) xor inputs(58) xor inputs(61) xor inputs(62) xor inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(191) <= inputs(250) xor inputs(251) xor inputs(254) xor inputs(255) ;
outputs(192) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(68) xor inputs(69) xor inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(87) xor inputs(88) xor inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(137) xor inputs(143) xor inputs(144) xor inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(193) <= inputs(64) xor inputs(65) xor inputs(68) xor inputs(69) xor inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(83) xor inputs(87) xor inputs(88) xor inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(136) xor inputs(137) xor inputs(143) xor inputs(144) xor inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(194) <= inputs(7) xor inputs(8) xor inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(136) xor inputs(137) xor inputs(143) xor inputs(144) xor inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(195) <= inputs(136) xor inputs(137) xor inputs(143) xor inputs(144) xor inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(196) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(6) xor inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(83) xor inputs(87) xor inputs(88) xor inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(197) <= inputs(83) xor inputs(87) xor inputs(88) xor inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(198) <= inputs(20) xor inputs(21) xor inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(199) <= inputs(198) xor inputs(199) xor inputs(206) xor inputs(207) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(200) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(68) xor inputs(69) xor inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(201) <= inputs(68) xor inputs(69) xor inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(202) <= inputs(8) xor inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(203) <= inputs(166) xor inputs(167) xor inputs(174) xor inputs(175) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(204) <= inputs(0) xor inputs(1) xor inputs(5) xor inputs(6) xor inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(205) <= inputs(109) xor inputs(110) xor inputs(117) xor inputs(118) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(206) <= inputs(37) xor inputs(38) xor inputs(45) xor inputs(46) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(207) <= inputs(230) xor inputs(231) xor inputs(238) xor inputs(239) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(208) <= inputs(1) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(209) <= inputs(64) xor inputs(65) xor inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(210) <= inputs(7) xor inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(211) <= inputs(150) xor inputs(151) xor inputs(158) xor inputs(159) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(212) <= inputs(1) xor inputs(5) xor inputs(6) xor inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(213) <= inputs(94) xor inputs(95) xor inputs(102) xor inputs(103) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(214) <= inputs(24) xor inputs(25) xor inputs(32) xor inputs(33) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(215) <= inputs(214) xor inputs(215) xor inputs(222) xor inputs(223) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(216) <= inputs(1) xor inputs(5) xor inputs(6) xor inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(217) <= inputs(73) xor inputs(74) xor inputs(81) xor inputs(82) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(218) <= inputs(10) xor inputs(11) xor inputs(17) xor inputs(18) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(219) <= inputs(182) xor inputs(183) xor inputs(190) xor inputs(191) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(220) <= inputs(1) xor inputs(5) xor inputs(6) xor inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(221) <= inputs(125) xor inputs(126) xor inputs(133) xor inputs(134) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(222) <= inputs(53) xor inputs(54) xor inputs(61) xor inputs(62) xor inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(223) <= inputs(246) xor inputs(247) xor inputs(254) xor inputs(255) ;
outputs(224) <= inputs(0) xor inputs(5) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(32) xor inputs(33) xor inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(68) xor inputs(69) xor inputs(81) xor inputs(82) xor inputs(87) xor inputs(88) xor inputs(102) xor inputs(103) xor inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(143) xor inputs(144) xor inputs(158) xor inputs(159) xor inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(225) <= inputs(64) xor inputs(65) xor inputs(68) xor inputs(69) xor inputs(81) xor inputs(82) xor inputs(87) xor inputs(88) xor inputs(102) xor inputs(103) xor inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(143) xor inputs(144) xor inputs(158) xor inputs(159) xor inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(226) <= inputs(7) xor inputs(8) xor inputs(17) xor inputs(18) xor inputs(20) xor inputs(21) xor inputs(32) xor inputs(33) xor inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(143) xor inputs(144) xor inputs(158) xor inputs(159) xor inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(227) <= inputs(143) xor inputs(144) xor inputs(158) xor inputs(159) xor inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(228) <= inputs(0) xor inputs(5) xor inputs(6) xor inputs(20) xor inputs(21) xor inputs(32) xor inputs(33) xor inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(87) xor inputs(88) xor inputs(102) xor inputs(103) xor inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(229) <= inputs(87) xor inputs(88) xor inputs(102) xor inputs(103) xor inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(230) <= inputs(20) xor inputs(21) xor inputs(32) xor inputs(33) xor inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(231) <= inputs(206) xor inputs(207) xor inputs(222) xor inputs(223) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(232) <= inputs(0) xor inputs(5) xor inputs(6) xor inputs(8) xor inputs(17) xor inputs(18) xor inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(68) xor inputs(69) xor inputs(81) xor inputs(82) xor inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(233) <= inputs(68) xor inputs(69) xor inputs(81) xor inputs(82) xor inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(234) <= inputs(8) xor inputs(17) xor inputs(18) xor inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(235) <= inputs(174) xor inputs(175) xor inputs(190) xor inputs(191) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(236) <= inputs(0) xor inputs(5) xor inputs(6) xor inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(237) <= inputs(117) xor inputs(118) xor inputs(133) xor inputs(134) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(238) <= inputs(45) xor inputs(46) xor inputs(61) xor inputs(62) xor inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(239) <= inputs(238) xor inputs(239) xor inputs(254) xor inputs(255) ;
outputs(240) <= inputs(5) xor inputs(6) xor inputs(7) xor inputs(17) xor inputs(18) xor inputs(32) xor inputs(33) xor inputs(61) xor inputs(62) xor inputs(64) xor inputs(65) xor inputs(81) xor inputs(82) xor inputs(102) xor inputs(103) xor inputs(133) xor inputs(134) xor inputs(158) xor inputs(159) xor inputs(190) xor inputs(191) xor inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(241) <= inputs(64) xor inputs(65) xor inputs(81) xor inputs(82) xor inputs(102) xor inputs(103) xor inputs(133) xor inputs(134) xor inputs(158) xor inputs(159) xor inputs(190) xor inputs(191) xor inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(242) <= inputs(7) xor inputs(17) xor inputs(18) xor inputs(32) xor inputs(33) xor inputs(61) xor inputs(62) xor inputs(158) xor inputs(159) xor inputs(190) xor inputs(191) xor inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(243) <= inputs(158) xor inputs(159) xor inputs(190) xor inputs(191) xor inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(244) <= inputs(5) xor inputs(6) xor inputs(32) xor inputs(33) xor inputs(61) xor inputs(62) xor inputs(102) xor inputs(103) xor inputs(133) xor inputs(134) xor inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(245) <= inputs(102) xor inputs(103) xor inputs(133) xor inputs(134) xor inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(246) <= inputs(32) xor inputs(33) xor inputs(61) xor inputs(62) xor inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(247) <= inputs(222) xor inputs(223) xor inputs(254) xor inputs(255) ;
outputs(248) <= inputs(5) xor inputs(6) xor inputs(17) xor inputs(18) xor inputs(61) xor inputs(62) xor inputs(81) xor inputs(82) xor inputs(133) xor inputs(134) xor inputs(190) xor inputs(191) xor inputs(254) xor inputs(255) ;
outputs(249) <= inputs(81) xor inputs(82) xor inputs(133) xor inputs(134) xor inputs(190) xor inputs(191) xor inputs(254) xor inputs(255) ;
outputs(250) <= inputs(17) xor inputs(18) xor inputs(61) xor inputs(62) xor inputs(190) xor inputs(191) xor inputs(254) xor inputs(255) ;
outputs(251) <= inputs(190) xor inputs(191) xor inputs(254) xor inputs(255) ;
outputs(252) <= inputs(5) xor inputs(6) xor inputs(61) xor inputs(62) xor inputs(133) xor inputs(134) xor inputs(254) xor inputs(255) ;
outputs(253) <= inputs(133) xor inputs(134) xor inputs(254) xor inputs(255) ;
outputs(254) <= inputs(61) xor inputs(62) xor inputs(254) xor inputs(255) ;
outputs(255) <= inputs(254) xor inputs(255) ;
outputs(256) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(135) xor inputs(137) xor inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(257) <= inputs(63) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(135) xor inputs(137) xor inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(258) <= inputs(7) xor inputs(8) xor inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(135) xor inputs(137) xor inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(259) <= inputs(135) xor inputs(137) xor inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(260) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(83) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(261) <= inputs(83) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(262) <= inputs(19) xor inputs(21) xor inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(263) <= inputs(193) xor inputs(195) xor inputs(197) xor inputs(199) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(264) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(8) xor inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(265) <= inputs(66) xor inputs(67) xor inputs(69) xor inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(266) <= inputs(8) xor inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(267) <= inputs(161) xor inputs(163) xor inputs(165) xor inputs(167) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(268) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(269) <= inputs(104) xor inputs(106) xor inputs(108) xor inputs(110) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(270) <= inputs(34) xor inputs(36) xor inputs(38) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(271) <= inputs(225) xor inputs(227) xor inputs(229) xor inputs(231) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(272) <= inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(273) <= inputs(63) xor inputs(65) xor inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(274) <= inputs(7) xor inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(275) <= inputs(145) xor inputs(147) xor inputs(149) xor inputs(151) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(276) <= inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(277) <= inputs(89) xor inputs(91) xor inputs(93) xor inputs(95) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(278) <= inputs(22) xor inputs(23) xor inputs(25) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(279) <= inputs(209) xor inputs(211) xor inputs(213) xor inputs(215) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(280) <= inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(281) <= inputs(70) xor inputs(72) xor inputs(74) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(282) <= inputs(9) xor inputs(11) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(283) <= inputs(177) xor inputs(179) xor inputs(181) xor inputs(183) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(284) <= inputs(1) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(285) <= inputs(120) xor inputs(122) xor inputs(124) xor inputs(126) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(286) <= inputs(48) xor inputs(50) xor inputs(52) xor inputs(54) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(287) <= inputs(241) xor inputs(243) xor inputs(245) xor inputs(247) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(288) <= inputs(0) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(289) <= inputs(63) xor inputs(65) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(290) <= inputs(7) xor inputs(8) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(291) <= inputs(138) xor inputs(140) xor inputs(142) xor inputs(144) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(292) <= inputs(0) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(19) xor inputs(21) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(84) xor inputs(86) xor inputs(88) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(293) <= inputs(84) xor inputs(86) xor inputs(88) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(294) <= inputs(19) xor inputs(21) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(295) <= inputs(201) xor inputs(203) xor inputs(205) xor inputs(207) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(296) <= inputs(0) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(8) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(66) xor inputs(67) xor inputs(69) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(297) <= inputs(66) xor inputs(67) xor inputs(69) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(298) <= inputs(8) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(299) <= inputs(169) xor inputs(171) xor inputs(173) xor inputs(175) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(300) <= inputs(0) xor inputs(2) xor inputs(4) xor inputs(6) xor inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(301) <= inputs(112) xor inputs(114) xor inputs(116) xor inputs(118) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(302) <= inputs(40) xor inputs(42) xor inputs(44) xor inputs(46) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(303) <= inputs(233) xor inputs(235) xor inputs(237) xor inputs(239) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(304) <= inputs(2) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(305) <= inputs(63) xor inputs(65) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(306) <= inputs(7) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(307) <= inputs(153) xor inputs(155) xor inputs(157) xor inputs(159) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(308) <= inputs(2) xor inputs(4) xor inputs(6) xor inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(309) <= inputs(97) xor inputs(99) xor inputs(101) xor inputs(103) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(310) <= inputs(27) xor inputs(29) xor inputs(31) xor inputs(33) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(311) <= inputs(217) xor inputs(219) xor inputs(221) xor inputs(223) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(312) <= inputs(2) xor inputs(4) xor inputs(6) xor inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(313) <= inputs(76) xor inputs(78) xor inputs(80) xor inputs(82) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(314) <= inputs(12) xor inputs(14) xor inputs(16) xor inputs(18) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(315) <= inputs(185) xor inputs(187) xor inputs(189) xor inputs(191) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(316) <= inputs(2) xor inputs(4) xor inputs(6) xor inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(317) <= inputs(128) xor inputs(130) xor inputs(132) xor inputs(134) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(318) <= inputs(56) xor inputs(58) xor inputs(60) xor inputs(62) xor inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(319) <= inputs(249) xor inputs(251) xor inputs(253) xor inputs(255) ;
outputs(320) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(83) xor inputs(86) xor inputs(88) xor inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(135) xor inputs(137) xor inputs(142) xor inputs(144) xor inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(321) <= inputs(63) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(83) xor inputs(86) xor inputs(88) xor inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(135) xor inputs(137) xor inputs(142) xor inputs(144) xor inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(322) <= inputs(7) xor inputs(8) xor inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(135) xor inputs(137) xor inputs(142) xor inputs(144) xor inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(323) <= inputs(135) xor inputs(137) xor inputs(142) xor inputs(144) xor inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(324) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(6) xor inputs(19) xor inputs(21) xor inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(83) xor inputs(86) xor inputs(88) xor inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(325) <= inputs(83) xor inputs(86) xor inputs(88) xor inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(326) <= inputs(19) xor inputs(21) xor inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(327) <= inputs(197) xor inputs(199) xor inputs(205) xor inputs(207) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(328) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(6) xor inputs(8) xor inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(67) xor inputs(69) xor inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(329) <= inputs(67) xor inputs(69) xor inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(330) <= inputs(8) xor inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(331) <= inputs(165) xor inputs(167) xor inputs(173) xor inputs(175) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(332) <= inputs(0) xor inputs(1) xor inputs(4) xor inputs(6) xor inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(333) <= inputs(108) xor inputs(110) xor inputs(116) xor inputs(118) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(334) <= inputs(36) xor inputs(38) xor inputs(44) xor inputs(46) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(335) <= inputs(229) xor inputs(231) xor inputs(237) xor inputs(239) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(336) <= inputs(1) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(337) <= inputs(63) xor inputs(65) xor inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(338) <= inputs(7) xor inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(339) <= inputs(149) xor inputs(151) xor inputs(157) xor inputs(159) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(340) <= inputs(1) xor inputs(4) xor inputs(6) xor inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(341) <= inputs(93) xor inputs(95) xor inputs(101) xor inputs(103) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(342) <= inputs(23) xor inputs(25) xor inputs(31) xor inputs(33) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(343) <= inputs(213) xor inputs(215) xor inputs(221) xor inputs(223) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(344) <= inputs(1) xor inputs(4) xor inputs(6) xor inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(345) <= inputs(72) xor inputs(74) xor inputs(80) xor inputs(82) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(346) <= inputs(9) xor inputs(11) xor inputs(16) xor inputs(18) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(347) <= inputs(181) xor inputs(183) xor inputs(189) xor inputs(191) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(348) <= inputs(1) xor inputs(4) xor inputs(6) xor inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(349) <= inputs(124) xor inputs(126) xor inputs(132) xor inputs(134) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(350) <= inputs(52) xor inputs(54) xor inputs(60) xor inputs(62) xor inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(351) <= inputs(245) xor inputs(247) xor inputs(253) xor inputs(255) ;
outputs(352) <= inputs(0) xor inputs(4) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(31) xor inputs(33) xor inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(80) xor inputs(82) xor inputs(86) xor inputs(88) xor inputs(101) xor inputs(103) xor inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(142) xor inputs(144) xor inputs(157) xor inputs(159) xor inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(353) <= inputs(63) xor inputs(65) xor inputs(67) xor inputs(69) xor inputs(80) xor inputs(82) xor inputs(86) xor inputs(88) xor inputs(101) xor inputs(103) xor inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(142) xor inputs(144) xor inputs(157) xor inputs(159) xor inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(354) <= inputs(7) xor inputs(8) xor inputs(16) xor inputs(18) xor inputs(19) xor inputs(21) xor inputs(31) xor inputs(33) xor inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(142) xor inputs(144) xor inputs(157) xor inputs(159) xor inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(355) <= inputs(142) xor inputs(144) xor inputs(157) xor inputs(159) xor inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(356) <= inputs(0) xor inputs(4) xor inputs(6) xor inputs(19) xor inputs(21) xor inputs(31) xor inputs(33) xor inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(86) xor inputs(88) xor inputs(101) xor inputs(103) xor inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(357) <= inputs(86) xor inputs(88) xor inputs(101) xor inputs(103) xor inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(358) <= inputs(19) xor inputs(21) xor inputs(31) xor inputs(33) xor inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(359) <= inputs(205) xor inputs(207) xor inputs(221) xor inputs(223) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(360) <= inputs(0) xor inputs(4) xor inputs(6) xor inputs(8) xor inputs(16) xor inputs(18) xor inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(67) xor inputs(69) xor inputs(80) xor inputs(82) xor inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(361) <= inputs(67) xor inputs(69) xor inputs(80) xor inputs(82) xor inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(362) <= inputs(8) xor inputs(16) xor inputs(18) xor inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(363) <= inputs(173) xor inputs(175) xor inputs(189) xor inputs(191) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(364) <= inputs(0) xor inputs(4) xor inputs(6) xor inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(365) <= inputs(116) xor inputs(118) xor inputs(132) xor inputs(134) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(366) <= inputs(44) xor inputs(46) xor inputs(60) xor inputs(62) xor inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(367) <= inputs(237) xor inputs(239) xor inputs(253) xor inputs(255) ;
outputs(368) <= inputs(4) xor inputs(6) xor inputs(7) xor inputs(16) xor inputs(18) xor inputs(31) xor inputs(33) xor inputs(60) xor inputs(62) xor inputs(63) xor inputs(65) xor inputs(80) xor inputs(82) xor inputs(101) xor inputs(103) xor inputs(132) xor inputs(134) xor inputs(157) xor inputs(159) xor inputs(189) xor inputs(191) xor inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(369) <= inputs(63) xor inputs(65) xor inputs(80) xor inputs(82) xor inputs(101) xor inputs(103) xor inputs(132) xor inputs(134) xor inputs(157) xor inputs(159) xor inputs(189) xor inputs(191) xor inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(370) <= inputs(7) xor inputs(16) xor inputs(18) xor inputs(31) xor inputs(33) xor inputs(60) xor inputs(62) xor inputs(157) xor inputs(159) xor inputs(189) xor inputs(191) xor inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(371) <= inputs(157) xor inputs(159) xor inputs(189) xor inputs(191) xor inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(372) <= inputs(4) xor inputs(6) xor inputs(31) xor inputs(33) xor inputs(60) xor inputs(62) xor inputs(101) xor inputs(103) xor inputs(132) xor inputs(134) xor inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(373) <= inputs(101) xor inputs(103) xor inputs(132) xor inputs(134) xor inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(374) <= inputs(31) xor inputs(33) xor inputs(60) xor inputs(62) xor inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(375) <= inputs(221) xor inputs(223) xor inputs(253) xor inputs(255) ;
outputs(376) <= inputs(4) xor inputs(6) xor inputs(16) xor inputs(18) xor inputs(60) xor inputs(62) xor inputs(80) xor inputs(82) xor inputs(132) xor inputs(134) xor inputs(189) xor inputs(191) xor inputs(253) xor inputs(255) ;
outputs(377) <= inputs(80) xor inputs(82) xor inputs(132) xor inputs(134) xor inputs(189) xor inputs(191) xor inputs(253) xor inputs(255) ;
outputs(378) <= inputs(16) xor inputs(18) xor inputs(60) xor inputs(62) xor inputs(189) xor inputs(191) xor inputs(253) xor inputs(255) ;
outputs(379) <= inputs(189) xor inputs(191) xor inputs(253) xor inputs(255) ;
outputs(380) <= inputs(4) xor inputs(6) xor inputs(60) xor inputs(62) xor inputs(132) xor inputs(134) xor inputs(253) xor inputs(255) ;
outputs(381) <= inputs(132) xor inputs(134) xor inputs(253) xor inputs(255) ;
outputs(382) <= inputs(60) xor inputs(62) xor inputs(253) xor inputs(255) ;
outputs(383) <= inputs(253) xor inputs(255) ;
outputs(384) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(11) xor inputs(14) xor inputs(18) xor inputs(21) xor inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(65) xor inputs(66) xor inputs(69) xor inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(88) xor inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(137) xor inputs(140) xor inputs(144) xor inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(385) <= inputs(65) xor inputs(66) xor inputs(69) xor inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(83) xor inputs(84) xor inputs(88) xor inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(137) xor inputs(140) xor inputs(144) xor inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(386) <= inputs(7) xor inputs(8) xor inputs(11) xor inputs(14) xor inputs(18) xor inputs(21) xor inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(137) xor inputs(140) xor inputs(144) xor inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(387) <= inputs(137) xor inputs(140) xor inputs(144) xor inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(388) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(6) xor inputs(21) xor inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(83) xor inputs(84) xor inputs(88) xor inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(389) <= inputs(83) xor inputs(84) xor inputs(88) xor inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(390) <= inputs(21) xor inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(391) <= inputs(195) xor inputs(199) xor inputs(203) xor inputs(207) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(392) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(6) xor inputs(8) xor inputs(11) xor inputs(14) xor inputs(18) xor inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(66) xor inputs(69) xor inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(393) <= inputs(66) xor inputs(69) xor inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(394) <= inputs(8) xor inputs(11) xor inputs(14) xor inputs(18) xor inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(395) <= inputs(163) xor inputs(167) xor inputs(171) xor inputs(175) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(396) <= inputs(0) xor inputs(1) xor inputs(2) xor inputs(6) xor inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(397) <= inputs(106) xor inputs(110) xor inputs(114) xor inputs(118) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(398) <= inputs(34) xor inputs(38) xor inputs(42) xor inputs(46) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(399) <= inputs(227) xor inputs(231) xor inputs(235) xor inputs(239) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(400) <= inputs(1) xor inputs(2) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(14) xor inputs(18) xor inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(65) xor inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(401) <= inputs(65) xor inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(402) <= inputs(7) xor inputs(11) xor inputs(14) xor inputs(18) xor inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(403) <= inputs(147) xor inputs(151) xor inputs(155) xor inputs(159) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(404) <= inputs(1) xor inputs(2) xor inputs(6) xor inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(405) <= inputs(91) xor inputs(95) xor inputs(99) xor inputs(103) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(406) <= inputs(22) xor inputs(25) xor inputs(29) xor inputs(33) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(407) <= inputs(211) xor inputs(215) xor inputs(219) xor inputs(223) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(408) <= inputs(1) xor inputs(2) xor inputs(6) xor inputs(11) xor inputs(14) xor inputs(18) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(409) <= inputs(70) xor inputs(74) xor inputs(78) xor inputs(82) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(410) <= inputs(11) xor inputs(14) xor inputs(18) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(411) <= inputs(179) xor inputs(183) xor inputs(187) xor inputs(191) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(412) <= inputs(1) xor inputs(2) xor inputs(6) xor inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(413) <= inputs(122) xor inputs(126) xor inputs(130) xor inputs(134) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(414) <= inputs(50) xor inputs(54) xor inputs(58) xor inputs(62) xor inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(415) <= inputs(243) xor inputs(247) xor inputs(251) xor inputs(255) ;
outputs(416) <= inputs(0) xor inputs(2) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(14) xor inputs(18) xor inputs(21) xor inputs(29) xor inputs(33) xor inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(65) xor inputs(66) xor inputs(69) xor inputs(78) xor inputs(82) xor inputs(84) xor inputs(88) xor inputs(99) xor inputs(103) xor inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(140) xor inputs(144) xor inputs(155) xor inputs(159) xor inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(417) <= inputs(65) xor inputs(66) xor inputs(69) xor inputs(78) xor inputs(82) xor inputs(84) xor inputs(88) xor inputs(99) xor inputs(103) xor inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(140) xor inputs(144) xor inputs(155) xor inputs(159) xor inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(418) <= inputs(7) xor inputs(8) xor inputs(14) xor inputs(18) xor inputs(21) xor inputs(29) xor inputs(33) xor inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(140) xor inputs(144) xor inputs(155) xor inputs(159) xor inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(419) <= inputs(140) xor inputs(144) xor inputs(155) xor inputs(159) xor inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(420) <= inputs(0) xor inputs(2) xor inputs(6) xor inputs(21) xor inputs(29) xor inputs(33) xor inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(84) xor inputs(88) xor inputs(99) xor inputs(103) xor inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(421) <= inputs(84) xor inputs(88) xor inputs(99) xor inputs(103) xor inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(422) <= inputs(21) xor inputs(29) xor inputs(33) xor inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(423) <= inputs(203) xor inputs(207) xor inputs(219) xor inputs(223) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(424) <= inputs(0) xor inputs(2) xor inputs(6) xor inputs(8) xor inputs(14) xor inputs(18) xor inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(66) xor inputs(69) xor inputs(78) xor inputs(82) xor inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(425) <= inputs(66) xor inputs(69) xor inputs(78) xor inputs(82) xor inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(426) <= inputs(8) xor inputs(14) xor inputs(18) xor inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(427) <= inputs(171) xor inputs(175) xor inputs(187) xor inputs(191) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(428) <= inputs(0) xor inputs(2) xor inputs(6) xor inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(429) <= inputs(114) xor inputs(118) xor inputs(130) xor inputs(134) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(430) <= inputs(42) xor inputs(46) xor inputs(58) xor inputs(62) xor inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(431) <= inputs(235) xor inputs(239) xor inputs(251) xor inputs(255) ;
outputs(432) <= inputs(2) xor inputs(6) xor inputs(7) xor inputs(14) xor inputs(18) xor inputs(29) xor inputs(33) xor inputs(58) xor inputs(62) xor inputs(65) xor inputs(78) xor inputs(82) xor inputs(99) xor inputs(103) xor inputs(130) xor inputs(134) xor inputs(155) xor inputs(159) xor inputs(187) xor inputs(191) xor inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(433) <= inputs(65) xor inputs(78) xor inputs(82) xor inputs(99) xor inputs(103) xor inputs(130) xor inputs(134) xor inputs(155) xor inputs(159) xor inputs(187) xor inputs(191) xor inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(434) <= inputs(7) xor inputs(14) xor inputs(18) xor inputs(29) xor inputs(33) xor inputs(58) xor inputs(62) xor inputs(155) xor inputs(159) xor inputs(187) xor inputs(191) xor inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(435) <= inputs(155) xor inputs(159) xor inputs(187) xor inputs(191) xor inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(436) <= inputs(2) xor inputs(6) xor inputs(29) xor inputs(33) xor inputs(58) xor inputs(62) xor inputs(99) xor inputs(103) xor inputs(130) xor inputs(134) xor inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(437) <= inputs(99) xor inputs(103) xor inputs(130) xor inputs(134) xor inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(438) <= inputs(29) xor inputs(33) xor inputs(58) xor inputs(62) xor inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(439) <= inputs(219) xor inputs(223) xor inputs(251) xor inputs(255) ;
outputs(440) <= inputs(2) xor inputs(6) xor inputs(14) xor inputs(18) xor inputs(58) xor inputs(62) xor inputs(78) xor inputs(82) xor inputs(130) xor inputs(134) xor inputs(187) xor inputs(191) xor inputs(251) xor inputs(255) ;
outputs(441) <= inputs(78) xor inputs(82) xor inputs(130) xor inputs(134) xor inputs(187) xor inputs(191) xor inputs(251) xor inputs(255) ;
outputs(442) <= inputs(14) xor inputs(18) xor inputs(58) xor inputs(62) xor inputs(187) xor inputs(191) xor inputs(251) xor inputs(255) ;
outputs(443) <= inputs(187) xor inputs(191) xor inputs(251) xor inputs(255) ;
outputs(444) <= inputs(2) xor inputs(6) xor inputs(58) xor inputs(62) xor inputs(130) xor inputs(134) xor inputs(251) xor inputs(255) ;
outputs(445) <= inputs(130) xor inputs(134) xor inputs(251) xor inputs(255) ;
outputs(446) <= inputs(58) xor inputs(62) xor inputs(251) xor inputs(255) ;
outputs(447) <= inputs(251) xor inputs(255) ;
outputs(448) <= inputs(0) xor inputs(1) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(11) xor inputs(18) xor inputs(21) xor inputs(25) xor inputs(33) xor inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(65) xor inputs(69) xor inputs(74) xor inputs(82) xor inputs(83) xor inputs(88) xor inputs(95) xor inputs(103) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(137) xor inputs(144) xor inputs(151) xor inputs(159) xor inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(449) <= inputs(65) xor inputs(69) xor inputs(74) xor inputs(82) xor inputs(83) xor inputs(88) xor inputs(95) xor inputs(103) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(137) xor inputs(144) xor inputs(151) xor inputs(159) xor inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(450) <= inputs(7) xor inputs(8) xor inputs(11) xor inputs(18) xor inputs(21) xor inputs(25) xor inputs(33) xor inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(137) xor inputs(144) xor inputs(151) xor inputs(159) xor inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(451) <= inputs(137) xor inputs(144) xor inputs(151) xor inputs(159) xor inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(452) <= inputs(0) xor inputs(1) xor inputs(6) xor inputs(21) xor inputs(25) xor inputs(33) xor inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(83) xor inputs(88) xor inputs(95) xor inputs(103) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(453) <= inputs(83) xor inputs(88) xor inputs(95) xor inputs(103) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(454) <= inputs(21) xor inputs(25) xor inputs(33) xor inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(455) <= inputs(199) xor inputs(207) xor inputs(215) xor inputs(223) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(456) <= inputs(0) xor inputs(1) xor inputs(6) xor inputs(8) xor inputs(11) xor inputs(18) xor inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(69) xor inputs(74) xor inputs(82) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(457) <= inputs(69) xor inputs(74) xor inputs(82) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(458) <= inputs(8) xor inputs(11) xor inputs(18) xor inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(459) <= inputs(167) xor inputs(175) xor inputs(183) xor inputs(191) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(460) <= inputs(0) xor inputs(1) xor inputs(6) xor inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(461) <= inputs(110) xor inputs(118) xor inputs(126) xor inputs(134) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(462) <= inputs(38) xor inputs(46) xor inputs(54) xor inputs(62) xor inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(463) <= inputs(231) xor inputs(239) xor inputs(247) xor inputs(255) ;
outputs(464) <= inputs(1) xor inputs(6) xor inputs(7) xor inputs(11) xor inputs(18) xor inputs(25) xor inputs(33) xor inputs(54) xor inputs(62) xor inputs(65) xor inputs(74) xor inputs(82) xor inputs(95) xor inputs(103) xor inputs(126) xor inputs(134) xor inputs(151) xor inputs(159) xor inputs(183) xor inputs(191) xor inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(465) <= inputs(65) xor inputs(74) xor inputs(82) xor inputs(95) xor inputs(103) xor inputs(126) xor inputs(134) xor inputs(151) xor inputs(159) xor inputs(183) xor inputs(191) xor inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(466) <= inputs(7) xor inputs(11) xor inputs(18) xor inputs(25) xor inputs(33) xor inputs(54) xor inputs(62) xor inputs(151) xor inputs(159) xor inputs(183) xor inputs(191) xor inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(467) <= inputs(151) xor inputs(159) xor inputs(183) xor inputs(191) xor inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(468) <= inputs(1) xor inputs(6) xor inputs(25) xor inputs(33) xor inputs(54) xor inputs(62) xor inputs(95) xor inputs(103) xor inputs(126) xor inputs(134) xor inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(469) <= inputs(95) xor inputs(103) xor inputs(126) xor inputs(134) xor inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(470) <= inputs(25) xor inputs(33) xor inputs(54) xor inputs(62) xor inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(471) <= inputs(215) xor inputs(223) xor inputs(247) xor inputs(255) ;
outputs(472) <= inputs(1) xor inputs(6) xor inputs(11) xor inputs(18) xor inputs(54) xor inputs(62) xor inputs(74) xor inputs(82) xor inputs(126) xor inputs(134) xor inputs(183) xor inputs(191) xor inputs(247) xor inputs(255) ;
outputs(473) <= inputs(74) xor inputs(82) xor inputs(126) xor inputs(134) xor inputs(183) xor inputs(191) xor inputs(247) xor inputs(255) ;
outputs(474) <= inputs(11) xor inputs(18) xor inputs(54) xor inputs(62) xor inputs(183) xor inputs(191) xor inputs(247) xor inputs(255) ;
outputs(475) <= inputs(183) xor inputs(191) xor inputs(247) xor inputs(255) ;
outputs(476) <= inputs(1) xor inputs(6) xor inputs(54) xor inputs(62) xor inputs(126) xor inputs(134) xor inputs(247) xor inputs(255) ;
outputs(477) <= inputs(126) xor inputs(134) xor inputs(247) xor inputs(255) ;
outputs(478) <= inputs(54) xor inputs(62) xor inputs(247) xor inputs(255) ;
outputs(479) <= inputs(247) xor inputs(255) ;
outputs(480) <= inputs(0) xor inputs(6) xor inputs(7) xor inputs(8) xor inputs(18) xor inputs(21) xor inputs(33) xor inputs(46) xor inputs(62) xor inputs(65) xor inputs(69) xor inputs(82) xor inputs(88) xor inputs(103) xor inputs(118) xor inputs(134) xor inputs(144) xor inputs(159) xor inputs(175) xor inputs(191) xor inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(481) <= inputs(65) xor inputs(69) xor inputs(82) xor inputs(88) xor inputs(103) xor inputs(118) xor inputs(134) xor inputs(144) xor inputs(159) xor inputs(175) xor inputs(191) xor inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(482) <= inputs(7) xor inputs(8) xor inputs(18) xor inputs(21) xor inputs(33) xor inputs(46) xor inputs(62) xor inputs(144) xor inputs(159) xor inputs(175) xor inputs(191) xor inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(483) <= inputs(144) xor inputs(159) xor inputs(175) xor inputs(191) xor inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(484) <= inputs(0) xor inputs(6) xor inputs(21) xor inputs(33) xor inputs(46) xor inputs(62) xor inputs(88) xor inputs(103) xor inputs(118) xor inputs(134) xor inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(485) <= inputs(88) xor inputs(103) xor inputs(118) xor inputs(134) xor inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(486) <= inputs(21) xor inputs(33) xor inputs(46) xor inputs(62) xor inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(487) <= inputs(207) xor inputs(223) xor inputs(239) xor inputs(255) ;
outputs(488) <= inputs(0) xor inputs(6) xor inputs(8) xor inputs(18) xor inputs(46) xor inputs(62) xor inputs(69) xor inputs(82) xor inputs(118) xor inputs(134) xor inputs(175) xor inputs(191) xor inputs(239) xor inputs(255) ;
outputs(489) <= inputs(69) xor inputs(82) xor inputs(118) xor inputs(134) xor inputs(175) xor inputs(191) xor inputs(239) xor inputs(255) ;
outputs(490) <= inputs(8) xor inputs(18) xor inputs(46) xor inputs(62) xor inputs(175) xor inputs(191) xor inputs(239) xor inputs(255) ;
outputs(491) <= inputs(175) xor inputs(191) xor inputs(239) xor inputs(255) ;
outputs(492) <= inputs(0) xor inputs(6) xor inputs(46) xor inputs(62) xor inputs(118) xor inputs(134) xor inputs(239) xor inputs(255) ;
outputs(493) <= inputs(118) xor inputs(134) xor inputs(239) xor inputs(255) ;
outputs(494) <= inputs(46) xor inputs(62) xor inputs(239) xor inputs(255) ;
outputs(495) <= inputs(239) xor inputs(255) ;
outputs(496) <= inputs(6) xor inputs(7) xor inputs(18) xor inputs(33) xor inputs(62) xor inputs(65) xor inputs(82) xor inputs(103) xor inputs(134) xor inputs(159) xor inputs(191) xor inputs(223) xor inputs(255) ;
outputs(497) <= inputs(65) xor inputs(82) xor inputs(103) xor inputs(134) xor inputs(159) xor inputs(191) xor inputs(223) xor inputs(255) ;
outputs(498) <= inputs(7) xor inputs(18) xor inputs(33) xor inputs(62) xor inputs(159) xor inputs(191) xor inputs(223) xor inputs(255) ;
outputs(499) <= inputs(159) xor inputs(191) xor inputs(223) xor inputs(255) ;
outputs(500) <= inputs(6) xor inputs(33) xor inputs(62) xor inputs(103) xor inputs(134) xor inputs(223) xor inputs(255) ;
outputs(501) <= inputs(103) xor inputs(134) xor inputs(223) xor inputs(255) ;
outputs(502) <= inputs(33) xor inputs(62) xor inputs(223) xor inputs(255) ;
outputs(503) <= inputs(223) xor inputs(255) ;
outputs(504) <= inputs(6) xor inputs(18) xor inputs(62) xor inputs(82) xor inputs(134) xor inputs(191) xor inputs(255) ;
outputs(505) <= inputs(82) xor inputs(134) xor inputs(191) xor inputs(255) ;
outputs(506) <= inputs(18) xor inputs(62) xor inputs(191) xor inputs(255) ;
outputs(507) <= inputs(191) xor inputs(255) ;
outputs(508) <= inputs(6) xor inputs(62) xor inputs(134) xor inputs(255) ;
outputs(509) <= inputs(134) xor inputs(255) ;
outputs(510) <= inputs(62) xor inputs(255) ;
outputs(511) <= inputs(255);

end Behavioral;
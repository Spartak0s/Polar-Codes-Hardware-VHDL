----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:10:49 02/17/2016 
-- Design Name: 
-- Module Name:    PartialSumGenerator - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.MyPackage.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PartialSumGenerator is
	Port (estimated : in std_logic_vector(N-2 downto 0);
			partial_sums : out s_2d);
end PartialSumGenerator;

architecture Behavioral of PartialSumGenerator is
	--gnal temp : s_2d;
begin
partial_sums(1)(0) <= estimated(0);
partial_sums(1)(1) <= estimated(512);
partial_sums(1)(2) <= estimated(256);
partial_sums(1)(3) <= estimated(768);
partial_sums(1)(4) <= estimated(128);
partial_sums(1)(5) <= estimated(640);
partial_sums(1)(6) <= estimated(384);
partial_sums(1)(7) <= estimated(896);
partial_sums(1)(8) <= estimated(64);
partial_sums(1)(9) <= estimated(576);
partial_sums(1)(10) <= estimated(320);
partial_sums(1)(11) <= estimated(832);
partial_sums(1)(12) <= estimated(192);
partial_sums(1)(13) <= estimated(704);
partial_sums(1)(14) <= estimated(448);
partial_sums(1)(15) <= estimated(960);
partial_sums(1)(16) <= estimated(32);
partial_sums(1)(17) <= estimated(544);
partial_sums(1)(18) <= estimated(288);
partial_sums(1)(19) <= estimated(800);
partial_sums(1)(20) <= estimated(160);
partial_sums(1)(21) <= estimated(672);
partial_sums(1)(22) <= estimated(416);
partial_sums(1)(23) <= estimated(928);
partial_sums(1)(24) <= estimated(96);
partial_sums(1)(25) <= estimated(608);
partial_sums(1)(26) <= estimated(352);
partial_sums(1)(27) <= estimated(864);
partial_sums(1)(28) <= estimated(224);
partial_sums(1)(29) <= estimated(736);
partial_sums(1)(30) <= estimated(480);
partial_sums(1)(31) <= estimated(992);
partial_sums(1)(32) <= estimated(16);
partial_sums(1)(33) <= estimated(528);
partial_sums(1)(34) <= estimated(272);
partial_sums(1)(35) <= estimated(784);
partial_sums(1)(36) <= estimated(144);
partial_sums(1)(37) <= estimated(656);
partial_sums(1)(38) <= estimated(400);
partial_sums(1)(39) <= estimated(912);
partial_sums(1)(40) <= estimated(80);
partial_sums(1)(41) <= estimated(592);
partial_sums(1)(42) <= estimated(336);
partial_sums(1)(43) <= estimated(848);
partial_sums(1)(44) <= estimated(208);
partial_sums(1)(45) <= estimated(720);
partial_sums(1)(46) <= estimated(464);
partial_sums(1)(47) <= estimated(976);
partial_sums(1)(48) <= estimated(48);
partial_sums(1)(49) <= estimated(560);
partial_sums(1)(50) <= estimated(304);
partial_sums(1)(51) <= estimated(816);
partial_sums(1)(52) <= estimated(176);
partial_sums(1)(53) <= estimated(688);
partial_sums(1)(54) <= estimated(432);
partial_sums(1)(55) <= estimated(944);
partial_sums(1)(56) <= estimated(112);
partial_sums(1)(57) <= estimated(624);
partial_sums(1)(58) <= estimated(368);
partial_sums(1)(59) <= estimated(880);
partial_sums(1)(60) <= estimated(240);
partial_sums(1)(61) <= estimated(752);
partial_sums(1)(62) <= estimated(496);
partial_sums(1)(63) <= estimated(1008);
partial_sums(1)(64) <= estimated(8);
partial_sums(1)(65) <= estimated(520);
partial_sums(1)(66) <= estimated(264);
partial_sums(1)(67) <= estimated(776);
partial_sums(1)(68) <= estimated(136);
partial_sums(1)(69) <= estimated(648);
partial_sums(1)(70) <= estimated(392);
partial_sums(1)(71) <= estimated(904);
partial_sums(1)(72) <= estimated(72);
partial_sums(1)(73) <= estimated(584);
partial_sums(1)(74) <= estimated(328);
partial_sums(1)(75) <= estimated(840);
partial_sums(1)(76) <= estimated(200);
partial_sums(1)(77) <= estimated(712);
partial_sums(1)(78) <= estimated(456);
partial_sums(1)(79) <= estimated(968);
partial_sums(1)(80) <= estimated(40);
partial_sums(1)(81) <= estimated(552);
partial_sums(1)(82) <= estimated(296);
partial_sums(1)(83) <= estimated(808);
partial_sums(1)(84) <= estimated(168);
partial_sums(1)(85) <= estimated(680);
partial_sums(1)(86) <= estimated(424);
partial_sums(1)(87) <= estimated(936);
partial_sums(1)(88) <= estimated(104);
partial_sums(1)(89) <= estimated(616);
partial_sums(1)(90) <= estimated(360);
partial_sums(1)(91) <= estimated(872);
partial_sums(1)(92) <= estimated(232);
partial_sums(1)(93) <= estimated(744);
partial_sums(1)(94) <= estimated(488);
partial_sums(1)(95) <= estimated(1000);
partial_sums(1)(96) <= estimated(24);
partial_sums(1)(97) <= estimated(536);
partial_sums(1)(98) <= estimated(280);
partial_sums(1)(99) <= estimated(792);
partial_sums(1)(100) <= estimated(152);
partial_sums(1)(101) <= estimated(664);
partial_sums(1)(102) <= estimated(408);
partial_sums(1)(103) <= estimated(920);
partial_sums(1)(104) <= estimated(88);
partial_sums(1)(105) <= estimated(600);
partial_sums(1)(106) <= estimated(344);
partial_sums(1)(107) <= estimated(856);
partial_sums(1)(108) <= estimated(216);
partial_sums(1)(109) <= estimated(728);
partial_sums(1)(110) <= estimated(472);
partial_sums(1)(111) <= estimated(984);
partial_sums(1)(112) <= estimated(56);
partial_sums(1)(113) <= estimated(568);
partial_sums(1)(114) <= estimated(312);
partial_sums(1)(115) <= estimated(824);
partial_sums(1)(116) <= estimated(184);
partial_sums(1)(117) <= estimated(696);
partial_sums(1)(118) <= estimated(440);
partial_sums(1)(119) <= estimated(952);
partial_sums(1)(120) <= estimated(120);
partial_sums(1)(121) <= estimated(632);
partial_sums(1)(122) <= estimated(376);
partial_sums(1)(123) <= estimated(888);
partial_sums(1)(124) <= estimated(248);
partial_sums(1)(125) <= estimated(760);
partial_sums(1)(126) <= estimated(504);
partial_sums(1)(127) <= estimated(1016);
partial_sums(1)(128) <= estimated(4);
partial_sums(1)(129) <= estimated(516);
partial_sums(1)(130) <= estimated(260);
partial_sums(1)(131) <= estimated(772);
partial_sums(1)(132) <= estimated(132);
partial_sums(1)(133) <= estimated(644);
partial_sums(1)(134) <= estimated(388);
partial_sums(1)(135) <= estimated(900);
partial_sums(1)(136) <= estimated(68);
partial_sums(1)(137) <= estimated(580);
partial_sums(1)(138) <= estimated(324);
partial_sums(1)(139) <= estimated(836);
partial_sums(1)(140) <= estimated(196);
partial_sums(1)(141) <= estimated(708);
partial_sums(1)(142) <= estimated(452);
partial_sums(1)(143) <= estimated(964);
partial_sums(1)(144) <= estimated(36);
partial_sums(1)(145) <= estimated(548);
partial_sums(1)(146) <= estimated(292);
partial_sums(1)(147) <= estimated(804);
partial_sums(1)(148) <= estimated(164);
partial_sums(1)(149) <= estimated(676);
partial_sums(1)(150) <= estimated(420);
partial_sums(1)(151) <= estimated(932);
partial_sums(1)(152) <= estimated(100);
partial_sums(1)(153) <= estimated(612);
partial_sums(1)(154) <= estimated(356);
partial_sums(1)(155) <= estimated(868);
partial_sums(1)(156) <= estimated(228);
partial_sums(1)(157) <= estimated(740);
partial_sums(1)(158) <= estimated(484);
partial_sums(1)(159) <= estimated(996);
partial_sums(1)(160) <= estimated(20);
partial_sums(1)(161) <= estimated(532);
partial_sums(1)(162) <= estimated(276);
partial_sums(1)(163) <= estimated(788);
partial_sums(1)(164) <= estimated(148);
partial_sums(1)(165) <= estimated(660);
partial_sums(1)(166) <= estimated(404);
partial_sums(1)(167) <= estimated(916);
partial_sums(1)(168) <= estimated(84);
partial_sums(1)(169) <= estimated(596);
partial_sums(1)(170) <= estimated(340);
partial_sums(1)(171) <= estimated(852);
partial_sums(1)(172) <= estimated(212);
partial_sums(1)(173) <= estimated(724);
partial_sums(1)(174) <= estimated(468);
partial_sums(1)(175) <= estimated(980);
partial_sums(1)(176) <= estimated(52);
partial_sums(1)(177) <= estimated(564);
partial_sums(1)(178) <= estimated(308);
partial_sums(1)(179) <= estimated(820);
partial_sums(1)(180) <= estimated(180);
partial_sums(1)(181) <= estimated(692);
partial_sums(1)(182) <= estimated(436);
partial_sums(1)(183) <= estimated(948);
partial_sums(1)(184) <= estimated(116);
partial_sums(1)(185) <= estimated(628);
partial_sums(1)(186) <= estimated(372);
partial_sums(1)(187) <= estimated(884);
partial_sums(1)(188) <= estimated(244);
partial_sums(1)(189) <= estimated(756);
partial_sums(1)(190) <= estimated(500);
partial_sums(1)(191) <= estimated(1012);
partial_sums(1)(192) <= estimated(12);
partial_sums(1)(193) <= estimated(524);
partial_sums(1)(194) <= estimated(268);
partial_sums(1)(195) <= estimated(780);
partial_sums(1)(196) <= estimated(140);
partial_sums(1)(197) <= estimated(652);
partial_sums(1)(198) <= estimated(396);
partial_sums(1)(199) <= estimated(908);
partial_sums(1)(200) <= estimated(76);
partial_sums(1)(201) <= estimated(588);
partial_sums(1)(202) <= estimated(332);
partial_sums(1)(203) <= estimated(844);
partial_sums(1)(204) <= estimated(204);
partial_sums(1)(205) <= estimated(716);
partial_sums(1)(206) <= estimated(460);
partial_sums(1)(207) <= estimated(972);
partial_sums(1)(208) <= estimated(44);
partial_sums(1)(209) <= estimated(556);
partial_sums(1)(210) <= estimated(300);
partial_sums(1)(211) <= estimated(812);
partial_sums(1)(212) <= estimated(172);
partial_sums(1)(213) <= estimated(684);
partial_sums(1)(214) <= estimated(428);
partial_sums(1)(215) <= estimated(940);
partial_sums(1)(216) <= estimated(108);
partial_sums(1)(217) <= estimated(620);
partial_sums(1)(218) <= estimated(364);
partial_sums(1)(219) <= estimated(876);
partial_sums(1)(220) <= estimated(236);
partial_sums(1)(221) <= estimated(748);
partial_sums(1)(222) <= estimated(492);
partial_sums(1)(223) <= estimated(1004);
partial_sums(1)(224) <= estimated(28);
partial_sums(1)(225) <= estimated(540);
partial_sums(1)(226) <= estimated(284);
partial_sums(1)(227) <= estimated(796);
partial_sums(1)(228) <= estimated(156);
partial_sums(1)(229) <= estimated(668);
partial_sums(1)(230) <= estimated(412);
partial_sums(1)(231) <= estimated(924);
partial_sums(1)(232) <= estimated(92);
partial_sums(1)(233) <= estimated(604);
partial_sums(1)(234) <= estimated(348);
partial_sums(1)(235) <= estimated(860);
partial_sums(1)(236) <= estimated(220);
partial_sums(1)(237) <= estimated(732);
partial_sums(1)(238) <= estimated(476);
partial_sums(1)(239) <= estimated(988);
partial_sums(1)(240) <= estimated(60);
partial_sums(1)(241) <= estimated(572);
partial_sums(1)(242) <= estimated(316);
partial_sums(1)(243) <= estimated(828);
partial_sums(1)(244) <= estimated(188);
partial_sums(1)(245) <= estimated(700);
partial_sums(1)(246) <= estimated(444);
partial_sums(1)(247) <= estimated(956);
partial_sums(1)(248) <= estimated(124);
partial_sums(1)(249) <= estimated(636);
partial_sums(1)(250) <= estimated(380);
partial_sums(1)(251) <= estimated(892);
partial_sums(1)(252) <= estimated(252);
partial_sums(1)(253) <= estimated(764);
partial_sums(1)(254) <= estimated(508);
partial_sums(1)(255) <= estimated(1020);
partial_sums(1)(256) <= estimated(2);
partial_sums(1)(257) <= estimated(514);
partial_sums(1)(258) <= estimated(258);
partial_sums(1)(259) <= estimated(770);
partial_sums(1)(260) <= estimated(130);
partial_sums(1)(261) <= estimated(642);
partial_sums(1)(262) <= estimated(386);
partial_sums(1)(263) <= estimated(898);
partial_sums(1)(264) <= estimated(66);
partial_sums(1)(265) <= estimated(578);
partial_sums(1)(266) <= estimated(322);
partial_sums(1)(267) <= estimated(834);
partial_sums(1)(268) <= estimated(194);
partial_sums(1)(269) <= estimated(706);
partial_sums(1)(270) <= estimated(450);
partial_sums(1)(271) <= estimated(962);
partial_sums(1)(272) <= estimated(34);
partial_sums(1)(273) <= estimated(546);
partial_sums(1)(274) <= estimated(290);
partial_sums(1)(275) <= estimated(802);
partial_sums(1)(276) <= estimated(162);
partial_sums(1)(277) <= estimated(674);
partial_sums(1)(278) <= estimated(418);
partial_sums(1)(279) <= estimated(930);
partial_sums(1)(280) <= estimated(98);
partial_sums(1)(281) <= estimated(610);
partial_sums(1)(282) <= estimated(354);
partial_sums(1)(283) <= estimated(866);
partial_sums(1)(284) <= estimated(226);
partial_sums(1)(285) <= estimated(738);
partial_sums(1)(286) <= estimated(482);
partial_sums(1)(287) <= estimated(994);
partial_sums(1)(288) <= estimated(18);
partial_sums(1)(289) <= estimated(530);
partial_sums(1)(290) <= estimated(274);
partial_sums(1)(291) <= estimated(786);
partial_sums(1)(292) <= estimated(146);
partial_sums(1)(293) <= estimated(658);
partial_sums(1)(294) <= estimated(402);
partial_sums(1)(295) <= estimated(914);
partial_sums(1)(296) <= estimated(82);
partial_sums(1)(297) <= estimated(594);
partial_sums(1)(298) <= estimated(338);
partial_sums(1)(299) <= estimated(850);
partial_sums(1)(300) <= estimated(210);
partial_sums(1)(301) <= estimated(722);
partial_sums(1)(302) <= estimated(466);
partial_sums(1)(303) <= estimated(978);
partial_sums(1)(304) <= estimated(50);
partial_sums(1)(305) <= estimated(562);
partial_sums(1)(306) <= estimated(306);
partial_sums(1)(307) <= estimated(818);
partial_sums(1)(308) <= estimated(178);
partial_sums(1)(309) <= estimated(690);
partial_sums(1)(310) <= estimated(434);
partial_sums(1)(311) <= estimated(946);
partial_sums(1)(312) <= estimated(114);
partial_sums(1)(313) <= estimated(626);
partial_sums(1)(314) <= estimated(370);
partial_sums(1)(315) <= estimated(882);
partial_sums(1)(316) <= estimated(242);
partial_sums(1)(317) <= estimated(754);
partial_sums(1)(318) <= estimated(498);
partial_sums(1)(319) <= estimated(1010);
partial_sums(1)(320) <= estimated(10);
partial_sums(1)(321) <= estimated(522);
partial_sums(1)(322) <= estimated(266);
partial_sums(1)(323) <= estimated(778);
partial_sums(1)(324) <= estimated(138);
partial_sums(1)(325) <= estimated(650);
partial_sums(1)(326) <= estimated(394);
partial_sums(1)(327) <= estimated(906);
partial_sums(1)(328) <= estimated(74);
partial_sums(1)(329) <= estimated(586);
partial_sums(1)(330) <= estimated(330);
partial_sums(1)(331) <= estimated(842);
partial_sums(1)(332) <= estimated(202);
partial_sums(1)(333) <= estimated(714);
partial_sums(1)(334) <= estimated(458);
partial_sums(1)(335) <= estimated(970);
partial_sums(1)(336) <= estimated(42);
partial_sums(1)(337) <= estimated(554);
partial_sums(1)(338) <= estimated(298);
partial_sums(1)(339) <= estimated(810);
partial_sums(1)(340) <= estimated(170);
partial_sums(1)(341) <= estimated(682);
partial_sums(1)(342) <= estimated(426);
partial_sums(1)(343) <= estimated(938);
partial_sums(1)(344) <= estimated(106);
partial_sums(1)(345) <= estimated(618);
partial_sums(1)(346) <= estimated(362);
partial_sums(1)(347) <= estimated(874);
partial_sums(1)(348) <= estimated(234);
partial_sums(1)(349) <= estimated(746);
partial_sums(1)(350) <= estimated(490);
partial_sums(1)(351) <= estimated(1002);
partial_sums(1)(352) <= estimated(26);
partial_sums(1)(353) <= estimated(538);
partial_sums(1)(354) <= estimated(282);
partial_sums(1)(355) <= estimated(794);
partial_sums(1)(356) <= estimated(154);
partial_sums(1)(357) <= estimated(666);
partial_sums(1)(358) <= estimated(410);
partial_sums(1)(359) <= estimated(922);
partial_sums(1)(360) <= estimated(90);
partial_sums(1)(361) <= estimated(602);
partial_sums(1)(362) <= estimated(346);
partial_sums(1)(363) <= estimated(858);
partial_sums(1)(364) <= estimated(218);
partial_sums(1)(365) <= estimated(730);
partial_sums(1)(366) <= estimated(474);
partial_sums(1)(367) <= estimated(986);
partial_sums(1)(368) <= estimated(58);
partial_sums(1)(369) <= estimated(570);
partial_sums(1)(370) <= estimated(314);
partial_sums(1)(371) <= estimated(826);
partial_sums(1)(372) <= estimated(186);
partial_sums(1)(373) <= estimated(698);
partial_sums(1)(374) <= estimated(442);
partial_sums(1)(375) <= estimated(954);
partial_sums(1)(376) <= estimated(122);
partial_sums(1)(377) <= estimated(634);
partial_sums(1)(378) <= estimated(378);
partial_sums(1)(379) <= estimated(890);
partial_sums(1)(380) <= estimated(250);
partial_sums(1)(381) <= estimated(762);
partial_sums(1)(382) <= estimated(506);
partial_sums(1)(383) <= estimated(1018);
partial_sums(1)(384) <= estimated(6);
partial_sums(1)(385) <= estimated(518);
partial_sums(1)(386) <= estimated(262);
partial_sums(1)(387) <= estimated(774);
partial_sums(1)(388) <= estimated(134);
partial_sums(1)(389) <= estimated(646);
partial_sums(1)(390) <= estimated(390);
partial_sums(1)(391) <= estimated(902);
partial_sums(1)(392) <= estimated(70);
partial_sums(1)(393) <= estimated(582);
partial_sums(1)(394) <= estimated(326);
partial_sums(1)(395) <= estimated(838);
partial_sums(1)(396) <= estimated(198);
partial_sums(1)(397) <= estimated(710);
partial_sums(1)(398) <= estimated(454);
partial_sums(1)(399) <= estimated(966);
partial_sums(1)(400) <= estimated(38);
partial_sums(1)(401) <= estimated(550);
partial_sums(1)(402) <= estimated(294);
partial_sums(1)(403) <= estimated(806);
partial_sums(1)(404) <= estimated(166);
partial_sums(1)(405) <= estimated(678);
partial_sums(1)(406) <= estimated(422);
partial_sums(1)(407) <= estimated(934);
partial_sums(1)(408) <= estimated(102);
partial_sums(1)(409) <= estimated(614);
partial_sums(1)(410) <= estimated(358);
partial_sums(1)(411) <= estimated(870);
partial_sums(1)(412) <= estimated(230);
partial_sums(1)(413) <= estimated(742);
partial_sums(1)(414) <= estimated(486);
partial_sums(1)(415) <= estimated(998);
partial_sums(1)(416) <= estimated(22);
partial_sums(1)(417) <= estimated(534);
partial_sums(1)(418) <= estimated(278);
partial_sums(1)(419) <= estimated(790);
partial_sums(1)(420) <= estimated(150);
partial_sums(1)(421) <= estimated(662);
partial_sums(1)(422) <= estimated(406);
partial_sums(1)(423) <= estimated(918);
partial_sums(1)(424) <= estimated(86);
partial_sums(1)(425) <= estimated(598);
partial_sums(1)(426) <= estimated(342);
partial_sums(1)(427) <= estimated(854);
partial_sums(1)(428) <= estimated(214);
partial_sums(1)(429) <= estimated(726);
partial_sums(1)(430) <= estimated(470);
partial_sums(1)(431) <= estimated(982);
partial_sums(1)(432) <= estimated(54);
partial_sums(1)(433) <= estimated(566);
partial_sums(1)(434) <= estimated(310);
partial_sums(1)(435) <= estimated(822);
partial_sums(1)(436) <= estimated(182);
partial_sums(1)(437) <= estimated(694);
partial_sums(1)(438) <= estimated(438);
partial_sums(1)(439) <= estimated(950);
partial_sums(1)(440) <= estimated(118);
partial_sums(1)(441) <= estimated(630);
partial_sums(1)(442) <= estimated(374);
partial_sums(1)(443) <= estimated(886);
partial_sums(1)(444) <= estimated(246);
partial_sums(1)(445) <= estimated(758);
partial_sums(1)(446) <= estimated(502);
partial_sums(1)(447) <= estimated(1014);
partial_sums(1)(448) <= estimated(14);
partial_sums(1)(449) <= estimated(526);
partial_sums(1)(450) <= estimated(270);
partial_sums(1)(451) <= estimated(782);
partial_sums(1)(452) <= estimated(142);
partial_sums(1)(453) <= estimated(654);
partial_sums(1)(454) <= estimated(398);
partial_sums(1)(455) <= estimated(910);
partial_sums(1)(456) <= estimated(78);
partial_sums(1)(457) <= estimated(590);
partial_sums(1)(458) <= estimated(334);
partial_sums(1)(459) <= estimated(846);
partial_sums(1)(460) <= estimated(206);
partial_sums(1)(461) <= estimated(718);
partial_sums(1)(462) <= estimated(462);
partial_sums(1)(463) <= estimated(974);
partial_sums(1)(464) <= estimated(46);
partial_sums(1)(465) <= estimated(558);
partial_sums(1)(466) <= estimated(302);
partial_sums(1)(467) <= estimated(814);
partial_sums(1)(468) <= estimated(174);
partial_sums(1)(469) <= estimated(686);
partial_sums(1)(470) <= estimated(430);
partial_sums(1)(471) <= estimated(942);
partial_sums(1)(472) <= estimated(110);
partial_sums(1)(473) <= estimated(622);
partial_sums(1)(474) <= estimated(366);
partial_sums(1)(475) <= estimated(878);
partial_sums(1)(476) <= estimated(238);
partial_sums(1)(477) <= estimated(750);
partial_sums(1)(478) <= estimated(494);
partial_sums(1)(479) <= estimated(1006);
partial_sums(1)(480) <= estimated(30);
partial_sums(1)(481) <= estimated(542);
partial_sums(1)(482) <= estimated(286);
partial_sums(1)(483) <= estimated(798);
partial_sums(1)(484) <= estimated(158);
partial_sums(1)(485) <= estimated(670);
partial_sums(1)(486) <= estimated(414);
partial_sums(1)(487) <= estimated(926);
partial_sums(1)(488) <= estimated(94);
partial_sums(1)(489) <= estimated(606);
partial_sums(1)(490) <= estimated(350);
partial_sums(1)(491) <= estimated(862);
partial_sums(1)(492) <= estimated(222);
partial_sums(1)(493) <= estimated(734);
partial_sums(1)(494) <= estimated(478);
partial_sums(1)(495) <= estimated(990);
partial_sums(1)(496) <= estimated(62);
partial_sums(1)(497) <= estimated(574);
partial_sums(1)(498) <= estimated(318);
partial_sums(1)(499) <= estimated(830);
partial_sums(1)(500) <= estimated(190);
partial_sums(1)(501) <= estimated(702);
partial_sums(1)(502) <= estimated(446);
partial_sums(1)(503) <= estimated(958);
partial_sums(1)(504) <= estimated(126);
partial_sums(1)(505) <= estimated(638);
partial_sums(1)(506) <= estimated(382);
partial_sums(1)(507) <= estimated(894);
partial_sums(1)(508) <= estimated(254);
partial_sums(1)(509) <= estimated(766);
partial_sums(1)(510) <= estimated(510);
partial_sums(1)(511) <= estimated(1022);
partial_sums(2)(0) <= estimated(0) xor estimated(1);
partial_sums(2)(1) <= estimated(512) xor estimated(513);
partial_sums(2)(2) <= estimated(256) xor estimated(257);
partial_sums(2)(3) <= estimated(768) xor estimated(769);
partial_sums(2)(4) <= estimated(128) xor estimated(129);
partial_sums(2)(5) <= estimated(640) xor estimated(641);
partial_sums(2)(6) <= estimated(384) xor estimated(385);
partial_sums(2)(7) <= estimated(896) xor estimated(897);
partial_sums(2)(8) <= estimated(64) xor estimated(65);
partial_sums(2)(9) <= estimated(576) xor estimated(577);
partial_sums(2)(10) <= estimated(320) xor estimated(321);
partial_sums(2)(11) <= estimated(832) xor estimated(833);
partial_sums(2)(12) <= estimated(192) xor estimated(193);
partial_sums(2)(13) <= estimated(704) xor estimated(705);
partial_sums(2)(14) <= estimated(448) xor estimated(449);
partial_sums(2)(15) <= estimated(960) xor estimated(961);
partial_sums(2)(16) <= estimated(32) xor estimated(33);
partial_sums(2)(17) <= estimated(544) xor estimated(545);
partial_sums(2)(18) <= estimated(288) xor estimated(289);
partial_sums(2)(19) <= estimated(800) xor estimated(801);
partial_sums(2)(20) <= estimated(160) xor estimated(161);
partial_sums(2)(21) <= estimated(672) xor estimated(673);
partial_sums(2)(22) <= estimated(416) xor estimated(417);
partial_sums(2)(23) <= estimated(928) xor estimated(929);
partial_sums(2)(24) <= estimated(96) xor estimated(97);
partial_sums(2)(25) <= estimated(608) xor estimated(609);
partial_sums(2)(26) <= estimated(352) xor estimated(353);
partial_sums(2)(27) <= estimated(864) xor estimated(865);
partial_sums(2)(28) <= estimated(224) xor estimated(225);
partial_sums(2)(29) <= estimated(736) xor estimated(737);
partial_sums(2)(30) <= estimated(480) xor estimated(481);
partial_sums(2)(31) <= estimated(992) xor estimated(993);
partial_sums(2)(32) <= estimated(16) xor estimated(17);
partial_sums(2)(33) <= estimated(528) xor estimated(529);
partial_sums(2)(34) <= estimated(272) xor estimated(273);
partial_sums(2)(35) <= estimated(784) xor estimated(785);
partial_sums(2)(36) <= estimated(144) xor estimated(145);
partial_sums(2)(37) <= estimated(656) xor estimated(657);
partial_sums(2)(38) <= estimated(400) xor estimated(401);
partial_sums(2)(39) <= estimated(912) xor estimated(913);
partial_sums(2)(40) <= estimated(80) xor estimated(81);
partial_sums(2)(41) <= estimated(592) xor estimated(593);
partial_sums(2)(42) <= estimated(336) xor estimated(337);
partial_sums(2)(43) <= estimated(848) xor estimated(849);
partial_sums(2)(44) <= estimated(208) xor estimated(209);
partial_sums(2)(45) <= estimated(720) xor estimated(721);
partial_sums(2)(46) <= estimated(464) xor estimated(465);
partial_sums(2)(47) <= estimated(976) xor estimated(977);
partial_sums(2)(48) <= estimated(48) xor estimated(49);
partial_sums(2)(49) <= estimated(560) xor estimated(561);
partial_sums(2)(50) <= estimated(304) xor estimated(305);
partial_sums(2)(51) <= estimated(816) xor estimated(817);
partial_sums(2)(52) <= estimated(176) xor estimated(177);
partial_sums(2)(53) <= estimated(688) xor estimated(689);
partial_sums(2)(54) <= estimated(432) xor estimated(433);
partial_sums(2)(55) <= estimated(944) xor estimated(945);
partial_sums(2)(56) <= estimated(112) xor estimated(113);
partial_sums(2)(57) <= estimated(624) xor estimated(625);
partial_sums(2)(58) <= estimated(368) xor estimated(369);
partial_sums(2)(59) <= estimated(880) xor estimated(881);
partial_sums(2)(60) <= estimated(240) xor estimated(241);
partial_sums(2)(61) <= estimated(752) xor estimated(753);
partial_sums(2)(62) <= estimated(496) xor estimated(497);
partial_sums(2)(63) <= estimated(1008) xor estimated(1009);
partial_sums(2)(64) <= estimated(8) xor estimated(9);
partial_sums(2)(65) <= estimated(520) xor estimated(521);
partial_sums(2)(66) <= estimated(264) xor estimated(265);
partial_sums(2)(67) <= estimated(776) xor estimated(777);
partial_sums(2)(68) <= estimated(136) xor estimated(137);
partial_sums(2)(69) <= estimated(648) xor estimated(649);
partial_sums(2)(70) <= estimated(392) xor estimated(393);
partial_sums(2)(71) <= estimated(904) xor estimated(905);
partial_sums(2)(72) <= estimated(72) xor estimated(73);
partial_sums(2)(73) <= estimated(584) xor estimated(585);
partial_sums(2)(74) <= estimated(328) xor estimated(329);
partial_sums(2)(75) <= estimated(840) xor estimated(841);
partial_sums(2)(76) <= estimated(200) xor estimated(201);
partial_sums(2)(77) <= estimated(712) xor estimated(713);
partial_sums(2)(78) <= estimated(456) xor estimated(457);
partial_sums(2)(79) <= estimated(968) xor estimated(969);
partial_sums(2)(80) <= estimated(40) xor estimated(41);
partial_sums(2)(81) <= estimated(552) xor estimated(553);
partial_sums(2)(82) <= estimated(296) xor estimated(297);
partial_sums(2)(83) <= estimated(808) xor estimated(809);
partial_sums(2)(84) <= estimated(168) xor estimated(169);
partial_sums(2)(85) <= estimated(680) xor estimated(681);
partial_sums(2)(86) <= estimated(424) xor estimated(425);
partial_sums(2)(87) <= estimated(936) xor estimated(937);
partial_sums(2)(88) <= estimated(104) xor estimated(105);
partial_sums(2)(89) <= estimated(616) xor estimated(617);
partial_sums(2)(90) <= estimated(360) xor estimated(361);
partial_sums(2)(91) <= estimated(872) xor estimated(873);
partial_sums(2)(92) <= estimated(232) xor estimated(233);
partial_sums(2)(93) <= estimated(744) xor estimated(745);
partial_sums(2)(94) <= estimated(488) xor estimated(489);
partial_sums(2)(95) <= estimated(1000) xor estimated(1001);
partial_sums(2)(96) <= estimated(24) xor estimated(25);
partial_sums(2)(97) <= estimated(536) xor estimated(537);
partial_sums(2)(98) <= estimated(280) xor estimated(281);
partial_sums(2)(99) <= estimated(792) xor estimated(793);
partial_sums(2)(100) <= estimated(152) xor estimated(153);
partial_sums(2)(101) <= estimated(664) xor estimated(665);
partial_sums(2)(102) <= estimated(408) xor estimated(409);
partial_sums(2)(103) <= estimated(920) xor estimated(921);
partial_sums(2)(104) <= estimated(88) xor estimated(89);
partial_sums(2)(105) <= estimated(600) xor estimated(601);
partial_sums(2)(106) <= estimated(344) xor estimated(345);
partial_sums(2)(107) <= estimated(856) xor estimated(857);
partial_sums(2)(108) <= estimated(216) xor estimated(217);
partial_sums(2)(109) <= estimated(728) xor estimated(729);
partial_sums(2)(110) <= estimated(472) xor estimated(473);
partial_sums(2)(111) <= estimated(984) xor estimated(985);
partial_sums(2)(112) <= estimated(56) xor estimated(57);
partial_sums(2)(113) <= estimated(568) xor estimated(569);
partial_sums(2)(114) <= estimated(312) xor estimated(313);
partial_sums(2)(115) <= estimated(824) xor estimated(825);
partial_sums(2)(116) <= estimated(184) xor estimated(185);
partial_sums(2)(117) <= estimated(696) xor estimated(697);
partial_sums(2)(118) <= estimated(440) xor estimated(441);
partial_sums(2)(119) <= estimated(952) xor estimated(953);
partial_sums(2)(120) <= estimated(120) xor estimated(121);
partial_sums(2)(121) <= estimated(632) xor estimated(633);
partial_sums(2)(122) <= estimated(376) xor estimated(377);
partial_sums(2)(123) <= estimated(888) xor estimated(889);
partial_sums(2)(124) <= estimated(248) xor estimated(249);
partial_sums(2)(125) <= estimated(760) xor estimated(761);
partial_sums(2)(126) <= estimated(504) xor estimated(505);
partial_sums(2)(127) <= estimated(1016) xor estimated(1017);
partial_sums(2)(128) <= estimated(4) xor estimated(5);
partial_sums(2)(129) <= estimated(516) xor estimated(517);
partial_sums(2)(130) <= estimated(260) xor estimated(261);
partial_sums(2)(131) <= estimated(772) xor estimated(773);
partial_sums(2)(132) <= estimated(132) xor estimated(133);
partial_sums(2)(133) <= estimated(644) xor estimated(645);
partial_sums(2)(134) <= estimated(388) xor estimated(389);
partial_sums(2)(135) <= estimated(900) xor estimated(901);
partial_sums(2)(136) <= estimated(68) xor estimated(69);
partial_sums(2)(137) <= estimated(580) xor estimated(581);
partial_sums(2)(138) <= estimated(324) xor estimated(325);
partial_sums(2)(139) <= estimated(836) xor estimated(837);
partial_sums(2)(140) <= estimated(196) xor estimated(197);
partial_sums(2)(141) <= estimated(708) xor estimated(709);
partial_sums(2)(142) <= estimated(452) xor estimated(453);
partial_sums(2)(143) <= estimated(964) xor estimated(965);
partial_sums(2)(144) <= estimated(36) xor estimated(37);
partial_sums(2)(145) <= estimated(548) xor estimated(549);
partial_sums(2)(146) <= estimated(292) xor estimated(293);
partial_sums(2)(147) <= estimated(804) xor estimated(805);
partial_sums(2)(148) <= estimated(164) xor estimated(165);
partial_sums(2)(149) <= estimated(676) xor estimated(677);
partial_sums(2)(150) <= estimated(420) xor estimated(421);
partial_sums(2)(151) <= estimated(932) xor estimated(933);
partial_sums(2)(152) <= estimated(100) xor estimated(101);
partial_sums(2)(153) <= estimated(612) xor estimated(613);
partial_sums(2)(154) <= estimated(356) xor estimated(357);
partial_sums(2)(155) <= estimated(868) xor estimated(869);
partial_sums(2)(156) <= estimated(228) xor estimated(229);
partial_sums(2)(157) <= estimated(740) xor estimated(741);
partial_sums(2)(158) <= estimated(484) xor estimated(485);
partial_sums(2)(159) <= estimated(996) xor estimated(997);
partial_sums(2)(160) <= estimated(20) xor estimated(21);
partial_sums(2)(161) <= estimated(532) xor estimated(533);
partial_sums(2)(162) <= estimated(276) xor estimated(277);
partial_sums(2)(163) <= estimated(788) xor estimated(789);
partial_sums(2)(164) <= estimated(148) xor estimated(149);
partial_sums(2)(165) <= estimated(660) xor estimated(661);
partial_sums(2)(166) <= estimated(404) xor estimated(405);
partial_sums(2)(167) <= estimated(916) xor estimated(917);
partial_sums(2)(168) <= estimated(84) xor estimated(85);
partial_sums(2)(169) <= estimated(596) xor estimated(597);
partial_sums(2)(170) <= estimated(340) xor estimated(341);
partial_sums(2)(171) <= estimated(852) xor estimated(853);
partial_sums(2)(172) <= estimated(212) xor estimated(213);
partial_sums(2)(173) <= estimated(724) xor estimated(725);
partial_sums(2)(174) <= estimated(468) xor estimated(469);
partial_sums(2)(175) <= estimated(980) xor estimated(981);
partial_sums(2)(176) <= estimated(52) xor estimated(53);
partial_sums(2)(177) <= estimated(564) xor estimated(565);
partial_sums(2)(178) <= estimated(308) xor estimated(309);
partial_sums(2)(179) <= estimated(820) xor estimated(821);
partial_sums(2)(180) <= estimated(180) xor estimated(181);
partial_sums(2)(181) <= estimated(692) xor estimated(693);
partial_sums(2)(182) <= estimated(436) xor estimated(437);
partial_sums(2)(183) <= estimated(948) xor estimated(949);
partial_sums(2)(184) <= estimated(116) xor estimated(117);
partial_sums(2)(185) <= estimated(628) xor estimated(629);
partial_sums(2)(186) <= estimated(372) xor estimated(373);
partial_sums(2)(187) <= estimated(884) xor estimated(885);
partial_sums(2)(188) <= estimated(244) xor estimated(245);
partial_sums(2)(189) <= estimated(756) xor estimated(757);
partial_sums(2)(190) <= estimated(500) xor estimated(501);
partial_sums(2)(191) <= estimated(1012) xor estimated(1013);
partial_sums(2)(192) <= estimated(12) xor estimated(13);
partial_sums(2)(193) <= estimated(524) xor estimated(525);
partial_sums(2)(194) <= estimated(268) xor estimated(269);
partial_sums(2)(195) <= estimated(780) xor estimated(781);
partial_sums(2)(196) <= estimated(140) xor estimated(141);
partial_sums(2)(197) <= estimated(652) xor estimated(653);
partial_sums(2)(198) <= estimated(396) xor estimated(397);
partial_sums(2)(199) <= estimated(908) xor estimated(909);
partial_sums(2)(200) <= estimated(76) xor estimated(77);
partial_sums(2)(201) <= estimated(588) xor estimated(589);
partial_sums(2)(202) <= estimated(332) xor estimated(333);
partial_sums(2)(203) <= estimated(844) xor estimated(845);
partial_sums(2)(204) <= estimated(204) xor estimated(205);
partial_sums(2)(205) <= estimated(716) xor estimated(717);
partial_sums(2)(206) <= estimated(460) xor estimated(461);
partial_sums(2)(207) <= estimated(972) xor estimated(973);
partial_sums(2)(208) <= estimated(44) xor estimated(45);
partial_sums(2)(209) <= estimated(556) xor estimated(557);
partial_sums(2)(210) <= estimated(300) xor estimated(301);
partial_sums(2)(211) <= estimated(812) xor estimated(813);
partial_sums(2)(212) <= estimated(172) xor estimated(173);
partial_sums(2)(213) <= estimated(684) xor estimated(685);
partial_sums(2)(214) <= estimated(428) xor estimated(429);
partial_sums(2)(215) <= estimated(940) xor estimated(941);
partial_sums(2)(216) <= estimated(108) xor estimated(109);
partial_sums(2)(217) <= estimated(620) xor estimated(621);
partial_sums(2)(218) <= estimated(364) xor estimated(365);
partial_sums(2)(219) <= estimated(876) xor estimated(877);
partial_sums(2)(220) <= estimated(236) xor estimated(237);
partial_sums(2)(221) <= estimated(748) xor estimated(749);
partial_sums(2)(222) <= estimated(492) xor estimated(493);
partial_sums(2)(223) <= estimated(1004) xor estimated(1005);
partial_sums(2)(224) <= estimated(28) xor estimated(29);
partial_sums(2)(225) <= estimated(540) xor estimated(541);
partial_sums(2)(226) <= estimated(284) xor estimated(285);
partial_sums(2)(227) <= estimated(796) xor estimated(797);
partial_sums(2)(228) <= estimated(156) xor estimated(157);
partial_sums(2)(229) <= estimated(668) xor estimated(669);
partial_sums(2)(230) <= estimated(412) xor estimated(413);
partial_sums(2)(231) <= estimated(924) xor estimated(925);
partial_sums(2)(232) <= estimated(92) xor estimated(93);
partial_sums(2)(233) <= estimated(604) xor estimated(605);
partial_sums(2)(234) <= estimated(348) xor estimated(349);
partial_sums(2)(235) <= estimated(860) xor estimated(861);
partial_sums(2)(236) <= estimated(220) xor estimated(221);
partial_sums(2)(237) <= estimated(732) xor estimated(733);
partial_sums(2)(238) <= estimated(476) xor estimated(477);
partial_sums(2)(239) <= estimated(988) xor estimated(989);
partial_sums(2)(240) <= estimated(60) xor estimated(61);
partial_sums(2)(241) <= estimated(572) xor estimated(573);
partial_sums(2)(242) <= estimated(316) xor estimated(317);
partial_sums(2)(243) <= estimated(828) xor estimated(829);
partial_sums(2)(244) <= estimated(188) xor estimated(189);
partial_sums(2)(245) <= estimated(700) xor estimated(701);
partial_sums(2)(246) <= estimated(444) xor estimated(445);
partial_sums(2)(247) <= estimated(956) xor estimated(957);
partial_sums(2)(248) <= estimated(124) xor estimated(125);
partial_sums(2)(249) <= estimated(636) xor estimated(637);
partial_sums(2)(250) <= estimated(380) xor estimated(381);
partial_sums(2)(251) <= estimated(892) xor estimated(893);
partial_sums(2)(252) <= estimated(252) xor estimated(253);
partial_sums(2)(253) <= estimated(764) xor estimated(765);
partial_sums(2)(254) <= estimated(508) xor estimated(509);
partial_sums(2)(255) <= estimated(1020) xor estimated(1021);
partial_sums(2)(256) <= estimated(1);
partial_sums(2)(257) <= estimated(513);
partial_sums(2)(258) <= estimated(257);
partial_sums(2)(259) <= estimated(769);
partial_sums(2)(260) <= estimated(129);
partial_sums(2)(261) <= estimated(641);
partial_sums(2)(262) <= estimated(385);
partial_sums(2)(263) <= estimated(897);
partial_sums(2)(264) <= estimated(65);
partial_sums(2)(265) <= estimated(577);
partial_sums(2)(266) <= estimated(321);
partial_sums(2)(267) <= estimated(833);
partial_sums(2)(268) <= estimated(193);
partial_sums(2)(269) <= estimated(705);
partial_sums(2)(270) <= estimated(449);
partial_sums(2)(271) <= estimated(961);
partial_sums(2)(272) <= estimated(33);
partial_sums(2)(273) <= estimated(545);
partial_sums(2)(274) <= estimated(289);
partial_sums(2)(275) <= estimated(801);
partial_sums(2)(276) <= estimated(161);
partial_sums(2)(277) <= estimated(673);
partial_sums(2)(278) <= estimated(417);
partial_sums(2)(279) <= estimated(929);
partial_sums(2)(280) <= estimated(97);
partial_sums(2)(281) <= estimated(609);
partial_sums(2)(282) <= estimated(353);
partial_sums(2)(283) <= estimated(865);
partial_sums(2)(284) <= estimated(225);
partial_sums(2)(285) <= estimated(737);
partial_sums(2)(286) <= estimated(481);
partial_sums(2)(287) <= estimated(993);
partial_sums(2)(288) <= estimated(17);
partial_sums(2)(289) <= estimated(529);
partial_sums(2)(290) <= estimated(273);
partial_sums(2)(291) <= estimated(785);
partial_sums(2)(292) <= estimated(145);
partial_sums(2)(293) <= estimated(657);
partial_sums(2)(294) <= estimated(401);
partial_sums(2)(295) <= estimated(913);
partial_sums(2)(296) <= estimated(81);
partial_sums(2)(297) <= estimated(593);
partial_sums(2)(298) <= estimated(337);
partial_sums(2)(299) <= estimated(849);
partial_sums(2)(300) <= estimated(209);
partial_sums(2)(301) <= estimated(721);
partial_sums(2)(302) <= estimated(465);
partial_sums(2)(303) <= estimated(977);
partial_sums(2)(304) <= estimated(49);
partial_sums(2)(305) <= estimated(561);
partial_sums(2)(306) <= estimated(305);
partial_sums(2)(307) <= estimated(817);
partial_sums(2)(308) <= estimated(177);
partial_sums(2)(309) <= estimated(689);
partial_sums(2)(310) <= estimated(433);
partial_sums(2)(311) <= estimated(945);
partial_sums(2)(312) <= estimated(113);
partial_sums(2)(313) <= estimated(625);
partial_sums(2)(314) <= estimated(369);
partial_sums(2)(315) <= estimated(881);
partial_sums(2)(316) <= estimated(241);
partial_sums(2)(317) <= estimated(753);
partial_sums(2)(318) <= estimated(497);
partial_sums(2)(319) <= estimated(1009);
partial_sums(2)(320) <= estimated(9);
partial_sums(2)(321) <= estimated(521);
partial_sums(2)(322) <= estimated(265);
partial_sums(2)(323) <= estimated(777);
partial_sums(2)(324) <= estimated(137);
partial_sums(2)(325) <= estimated(649);
partial_sums(2)(326) <= estimated(393);
partial_sums(2)(327) <= estimated(905);
partial_sums(2)(328) <= estimated(73);
partial_sums(2)(329) <= estimated(585);
partial_sums(2)(330) <= estimated(329);
partial_sums(2)(331) <= estimated(841);
partial_sums(2)(332) <= estimated(201);
partial_sums(2)(333) <= estimated(713);
partial_sums(2)(334) <= estimated(457);
partial_sums(2)(335) <= estimated(969);
partial_sums(2)(336) <= estimated(41);
partial_sums(2)(337) <= estimated(553);
partial_sums(2)(338) <= estimated(297);
partial_sums(2)(339) <= estimated(809);
partial_sums(2)(340) <= estimated(169);
partial_sums(2)(341) <= estimated(681);
partial_sums(2)(342) <= estimated(425);
partial_sums(2)(343) <= estimated(937);
partial_sums(2)(344) <= estimated(105);
partial_sums(2)(345) <= estimated(617);
partial_sums(2)(346) <= estimated(361);
partial_sums(2)(347) <= estimated(873);
partial_sums(2)(348) <= estimated(233);
partial_sums(2)(349) <= estimated(745);
partial_sums(2)(350) <= estimated(489);
partial_sums(2)(351) <= estimated(1001);
partial_sums(2)(352) <= estimated(25);
partial_sums(2)(353) <= estimated(537);
partial_sums(2)(354) <= estimated(281);
partial_sums(2)(355) <= estimated(793);
partial_sums(2)(356) <= estimated(153);
partial_sums(2)(357) <= estimated(665);
partial_sums(2)(358) <= estimated(409);
partial_sums(2)(359) <= estimated(921);
partial_sums(2)(360) <= estimated(89);
partial_sums(2)(361) <= estimated(601);
partial_sums(2)(362) <= estimated(345);
partial_sums(2)(363) <= estimated(857);
partial_sums(2)(364) <= estimated(217);
partial_sums(2)(365) <= estimated(729);
partial_sums(2)(366) <= estimated(473);
partial_sums(2)(367) <= estimated(985);
partial_sums(2)(368) <= estimated(57);
partial_sums(2)(369) <= estimated(569);
partial_sums(2)(370) <= estimated(313);
partial_sums(2)(371) <= estimated(825);
partial_sums(2)(372) <= estimated(185);
partial_sums(2)(373) <= estimated(697);
partial_sums(2)(374) <= estimated(441);
partial_sums(2)(375) <= estimated(953);
partial_sums(2)(376) <= estimated(121);
partial_sums(2)(377) <= estimated(633);
partial_sums(2)(378) <= estimated(377);
partial_sums(2)(379) <= estimated(889);
partial_sums(2)(380) <= estimated(249);
partial_sums(2)(381) <= estimated(761);
partial_sums(2)(382) <= estimated(505);
partial_sums(2)(383) <= estimated(1017);
partial_sums(2)(384) <= estimated(5);
partial_sums(2)(385) <= estimated(517);
partial_sums(2)(386) <= estimated(261);
partial_sums(2)(387) <= estimated(773);
partial_sums(2)(388) <= estimated(133);
partial_sums(2)(389) <= estimated(645);
partial_sums(2)(390) <= estimated(389);
partial_sums(2)(391) <= estimated(901);
partial_sums(2)(392) <= estimated(69);
partial_sums(2)(393) <= estimated(581);
partial_sums(2)(394) <= estimated(325);
partial_sums(2)(395) <= estimated(837);
partial_sums(2)(396) <= estimated(197);
partial_sums(2)(397) <= estimated(709);
partial_sums(2)(398) <= estimated(453);
partial_sums(2)(399) <= estimated(965);
partial_sums(2)(400) <= estimated(37);
partial_sums(2)(401) <= estimated(549);
partial_sums(2)(402) <= estimated(293);
partial_sums(2)(403) <= estimated(805);
partial_sums(2)(404) <= estimated(165);
partial_sums(2)(405) <= estimated(677);
partial_sums(2)(406) <= estimated(421);
partial_sums(2)(407) <= estimated(933);
partial_sums(2)(408) <= estimated(101);
partial_sums(2)(409) <= estimated(613);
partial_sums(2)(410) <= estimated(357);
partial_sums(2)(411) <= estimated(869);
partial_sums(2)(412) <= estimated(229);
partial_sums(2)(413) <= estimated(741);
partial_sums(2)(414) <= estimated(485);
partial_sums(2)(415) <= estimated(997);
partial_sums(2)(416) <= estimated(21);
partial_sums(2)(417) <= estimated(533);
partial_sums(2)(418) <= estimated(277);
partial_sums(2)(419) <= estimated(789);
partial_sums(2)(420) <= estimated(149);
partial_sums(2)(421) <= estimated(661);
partial_sums(2)(422) <= estimated(405);
partial_sums(2)(423) <= estimated(917);
partial_sums(2)(424) <= estimated(85);
partial_sums(2)(425) <= estimated(597);
partial_sums(2)(426) <= estimated(341);
partial_sums(2)(427) <= estimated(853);
partial_sums(2)(428) <= estimated(213);
partial_sums(2)(429) <= estimated(725);
partial_sums(2)(430) <= estimated(469);
partial_sums(2)(431) <= estimated(981);
partial_sums(2)(432) <= estimated(53);
partial_sums(2)(433) <= estimated(565);
partial_sums(2)(434) <= estimated(309);
partial_sums(2)(435) <= estimated(821);
partial_sums(2)(436) <= estimated(181);
partial_sums(2)(437) <= estimated(693);
partial_sums(2)(438) <= estimated(437);
partial_sums(2)(439) <= estimated(949);
partial_sums(2)(440) <= estimated(117);
partial_sums(2)(441) <= estimated(629);
partial_sums(2)(442) <= estimated(373);
partial_sums(2)(443) <= estimated(885);
partial_sums(2)(444) <= estimated(245);
partial_sums(2)(445) <= estimated(757);
partial_sums(2)(446) <= estimated(501);
partial_sums(2)(447) <= estimated(1013);
partial_sums(2)(448) <= estimated(13);
partial_sums(2)(449) <= estimated(525);
partial_sums(2)(450) <= estimated(269);
partial_sums(2)(451) <= estimated(781);
partial_sums(2)(452) <= estimated(141);
partial_sums(2)(453) <= estimated(653);
partial_sums(2)(454) <= estimated(397);
partial_sums(2)(455) <= estimated(909);
partial_sums(2)(456) <= estimated(77);
partial_sums(2)(457) <= estimated(589);
partial_sums(2)(458) <= estimated(333);
partial_sums(2)(459) <= estimated(845);
partial_sums(2)(460) <= estimated(205);
partial_sums(2)(461) <= estimated(717);
partial_sums(2)(462) <= estimated(461);
partial_sums(2)(463) <= estimated(973);
partial_sums(2)(464) <= estimated(45);
partial_sums(2)(465) <= estimated(557);
partial_sums(2)(466) <= estimated(301);
partial_sums(2)(467) <= estimated(813);
partial_sums(2)(468) <= estimated(173);
partial_sums(2)(469) <= estimated(685);
partial_sums(2)(470) <= estimated(429);
partial_sums(2)(471) <= estimated(941);
partial_sums(2)(472) <= estimated(109);
partial_sums(2)(473) <= estimated(621);
partial_sums(2)(474) <= estimated(365);
partial_sums(2)(475) <= estimated(877);
partial_sums(2)(476) <= estimated(237);
partial_sums(2)(477) <= estimated(749);
partial_sums(2)(478) <= estimated(493);
partial_sums(2)(479) <= estimated(1005);
partial_sums(2)(480) <= estimated(29);
partial_sums(2)(481) <= estimated(541);
partial_sums(2)(482) <= estimated(285);
partial_sums(2)(483) <= estimated(797);
partial_sums(2)(484) <= estimated(157);
partial_sums(2)(485) <= estimated(669);
partial_sums(2)(486) <= estimated(413);
partial_sums(2)(487) <= estimated(925);
partial_sums(2)(488) <= estimated(93);
partial_sums(2)(489) <= estimated(605);
partial_sums(2)(490) <= estimated(349);
partial_sums(2)(491) <= estimated(861);
partial_sums(2)(492) <= estimated(221);
partial_sums(2)(493) <= estimated(733);
partial_sums(2)(494) <= estimated(477);
partial_sums(2)(495) <= estimated(989);
partial_sums(2)(496) <= estimated(61);
partial_sums(2)(497) <= estimated(573);
partial_sums(2)(498) <= estimated(317);
partial_sums(2)(499) <= estimated(829);
partial_sums(2)(500) <= estimated(189);
partial_sums(2)(501) <= estimated(701);
partial_sums(2)(502) <= estimated(445);
partial_sums(2)(503) <= estimated(957);
partial_sums(2)(504) <= estimated(125);
partial_sums(2)(505) <= estimated(637);
partial_sums(2)(506) <= estimated(381);
partial_sums(2)(507) <= estimated(893);
partial_sums(2)(508) <= estimated(253);
partial_sums(2)(509) <= estimated(765);
partial_sums(2)(510) <= estimated(509);
partial_sums(2)(511) <= estimated(1021);
partial_sums(3)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3);
partial_sums(3)(1) <= estimated(512) xor estimated(513) xor estimated(514) xor estimated(515);
partial_sums(3)(2) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259);
partial_sums(3)(3) <= estimated(768) xor estimated(769) xor estimated(770) xor estimated(771);
partial_sums(3)(4) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131);
partial_sums(3)(5) <= estimated(640) xor estimated(641) xor estimated(642) xor estimated(643);
partial_sums(3)(6) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387);
partial_sums(3)(7) <= estimated(896) xor estimated(897) xor estimated(898) xor estimated(899);
partial_sums(3)(8) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67);
partial_sums(3)(9) <= estimated(576) xor estimated(577) xor estimated(578) xor estimated(579);
partial_sums(3)(10) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323);
partial_sums(3)(11) <= estimated(832) xor estimated(833) xor estimated(834) xor estimated(835);
partial_sums(3)(12) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195);
partial_sums(3)(13) <= estimated(704) xor estimated(705) xor estimated(706) xor estimated(707);
partial_sums(3)(14) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451);
partial_sums(3)(15) <= estimated(960) xor estimated(961) xor estimated(962) xor estimated(963);
partial_sums(3)(16) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35);
partial_sums(3)(17) <= estimated(544) xor estimated(545) xor estimated(546) xor estimated(547);
partial_sums(3)(18) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291);
partial_sums(3)(19) <= estimated(800) xor estimated(801) xor estimated(802) xor estimated(803);
partial_sums(3)(20) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163);
partial_sums(3)(21) <= estimated(672) xor estimated(673) xor estimated(674) xor estimated(675);
partial_sums(3)(22) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419);
partial_sums(3)(23) <= estimated(928) xor estimated(929) xor estimated(930) xor estimated(931);
partial_sums(3)(24) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99);
partial_sums(3)(25) <= estimated(608) xor estimated(609) xor estimated(610) xor estimated(611);
partial_sums(3)(26) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355);
partial_sums(3)(27) <= estimated(864) xor estimated(865) xor estimated(866) xor estimated(867);
partial_sums(3)(28) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227);
partial_sums(3)(29) <= estimated(736) xor estimated(737) xor estimated(738) xor estimated(739);
partial_sums(3)(30) <= estimated(480) xor estimated(481) xor estimated(482) xor estimated(483);
partial_sums(3)(31) <= estimated(992) xor estimated(993) xor estimated(994) xor estimated(995);
partial_sums(3)(32) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19);
partial_sums(3)(33) <= estimated(528) xor estimated(529) xor estimated(530) xor estimated(531);
partial_sums(3)(34) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275);
partial_sums(3)(35) <= estimated(784) xor estimated(785) xor estimated(786) xor estimated(787);
partial_sums(3)(36) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147);
partial_sums(3)(37) <= estimated(656) xor estimated(657) xor estimated(658) xor estimated(659);
partial_sums(3)(38) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403);
partial_sums(3)(39) <= estimated(912) xor estimated(913) xor estimated(914) xor estimated(915);
partial_sums(3)(40) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83);
partial_sums(3)(41) <= estimated(592) xor estimated(593) xor estimated(594) xor estimated(595);
partial_sums(3)(42) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339);
partial_sums(3)(43) <= estimated(848) xor estimated(849) xor estimated(850) xor estimated(851);
partial_sums(3)(44) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211);
partial_sums(3)(45) <= estimated(720) xor estimated(721) xor estimated(722) xor estimated(723);
partial_sums(3)(46) <= estimated(464) xor estimated(465) xor estimated(466) xor estimated(467);
partial_sums(3)(47) <= estimated(976) xor estimated(977) xor estimated(978) xor estimated(979);
partial_sums(3)(48) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51);
partial_sums(3)(49) <= estimated(560) xor estimated(561) xor estimated(562) xor estimated(563);
partial_sums(3)(50) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307);
partial_sums(3)(51) <= estimated(816) xor estimated(817) xor estimated(818) xor estimated(819);
partial_sums(3)(52) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179);
partial_sums(3)(53) <= estimated(688) xor estimated(689) xor estimated(690) xor estimated(691);
partial_sums(3)(54) <= estimated(432) xor estimated(433) xor estimated(434) xor estimated(435);
partial_sums(3)(55) <= estimated(944) xor estimated(945) xor estimated(946) xor estimated(947);
partial_sums(3)(56) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115);
partial_sums(3)(57) <= estimated(624) xor estimated(625) xor estimated(626) xor estimated(627);
partial_sums(3)(58) <= estimated(368) xor estimated(369) xor estimated(370) xor estimated(371);
partial_sums(3)(59) <= estimated(880) xor estimated(881) xor estimated(882) xor estimated(883);
partial_sums(3)(60) <= estimated(240) xor estimated(241) xor estimated(242) xor estimated(243);
partial_sums(3)(61) <= estimated(752) xor estimated(753) xor estimated(754) xor estimated(755);
partial_sums(3)(62) <= estimated(496) xor estimated(497) xor estimated(498) xor estimated(499);
partial_sums(3)(63) <= estimated(1008) xor estimated(1009) xor estimated(1010) xor estimated(1011);
partial_sums(3)(64) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11);
partial_sums(3)(65) <= estimated(520) xor estimated(521) xor estimated(522) xor estimated(523);
partial_sums(3)(66) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267);
partial_sums(3)(67) <= estimated(776) xor estimated(777) xor estimated(778) xor estimated(779);
partial_sums(3)(68) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139);
partial_sums(3)(69) <= estimated(648) xor estimated(649) xor estimated(650) xor estimated(651);
partial_sums(3)(70) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395);
partial_sums(3)(71) <= estimated(904) xor estimated(905) xor estimated(906) xor estimated(907);
partial_sums(3)(72) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75);
partial_sums(3)(73) <= estimated(584) xor estimated(585) xor estimated(586) xor estimated(587);
partial_sums(3)(74) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331);
partial_sums(3)(75) <= estimated(840) xor estimated(841) xor estimated(842) xor estimated(843);
partial_sums(3)(76) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203);
partial_sums(3)(77) <= estimated(712) xor estimated(713) xor estimated(714) xor estimated(715);
partial_sums(3)(78) <= estimated(456) xor estimated(457) xor estimated(458) xor estimated(459);
partial_sums(3)(79) <= estimated(968) xor estimated(969) xor estimated(970) xor estimated(971);
partial_sums(3)(80) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43);
partial_sums(3)(81) <= estimated(552) xor estimated(553) xor estimated(554) xor estimated(555);
partial_sums(3)(82) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299);
partial_sums(3)(83) <= estimated(808) xor estimated(809) xor estimated(810) xor estimated(811);
partial_sums(3)(84) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171);
partial_sums(3)(85) <= estimated(680) xor estimated(681) xor estimated(682) xor estimated(683);
partial_sums(3)(86) <= estimated(424) xor estimated(425) xor estimated(426) xor estimated(427);
partial_sums(3)(87) <= estimated(936) xor estimated(937) xor estimated(938) xor estimated(939);
partial_sums(3)(88) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107);
partial_sums(3)(89) <= estimated(616) xor estimated(617) xor estimated(618) xor estimated(619);
partial_sums(3)(90) <= estimated(360) xor estimated(361) xor estimated(362) xor estimated(363);
partial_sums(3)(91) <= estimated(872) xor estimated(873) xor estimated(874) xor estimated(875);
partial_sums(3)(92) <= estimated(232) xor estimated(233) xor estimated(234) xor estimated(235);
partial_sums(3)(93) <= estimated(744) xor estimated(745) xor estimated(746) xor estimated(747);
partial_sums(3)(94) <= estimated(488) xor estimated(489) xor estimated(490) xor estimated(491);
partial_sums(3)(95) <= estimated(1000) xor estimated(1001) xor estimated(1002) xor estimated(1003);
partial_sums(3)(96) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27);
partial_sums(3)(97) <= estimated(536) xor estimated(537) xor estimated(538) xor estimated(539);
partial_sums(3)(98) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283);
partial_sums(3)(99) <= estimated(792) xor estimated(793) xor estimated(794) xor estimated(795);
partial_sums(3)(100) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155);
partial_sums(3)(101) <= estimated(664) xor estimated(665) xor estimated(666) xor estimated(667);
partial_sums(3)(102) <= estimated(408) xor estimated(409) xor estimated(410) xor estimated(411);
partial_sums(3)(103) <= estimated(920) xor estimated(921) xor estimated(922) xor estimated(923);
partial_sums(3)(104) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91);
partial_sums(3)(105) <= estimated(600) xor estimated(601) xor estimated(602) xor estimated(603);
partial_sums(3)(106) <= estimated(344) xor estimated(345) xor estimated(346) xor estimated(347);
partial_sums(3)(107) <= estimated(856) xor estimated(857) xor estimated(858) xor estimated(859);
partial_sums(3)(108) <= estimated(216) xor estimated(217) xor estimated(218) xor estimated(219);
partial_sums(3)(109) <= estimated(728) xor estimated(729) xor estimated(730) xor estimated(731);
partial_sums(3)(110) <= estimated(472) xor estimated(473) xor estimated(474) xor estimated(475);
partial_sums(3)(111) <= estimated(984) xor estimated(985) xor estimated(986) xor estimated(987);
partial_sums(3)(112) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59);
partial_sums(3)(113) <= estimated(568) xor estimated(569) xor estimated(570) xor estimated(571);
partial_sums(3)(114) <= estimated(312) xor estimated(313) xor estimated(314) xor estimated(315);
partial_sums(3)(115) <= estimated(824) xor estimated(825) xor estimated(826) xor estimated(827);
partial_sums(3)(116) <= estimated(184) xor estimated(185) xor estimated(186) xor estimated(187);
partial_sums(3)(117) <= estimated(696) xor estimated(697) xor estimated(698) xor estimated(699);
partial_sums(3)(118) <= estimated(440) xor estimated(441) xor estimated(442) xor estimated(443);
partial_sums(3)(119) <= estimated(952) xor estimated(953) xor estimated(954) xor estimated(955);
partial_sums(3)(120) <= estimated(120) xor estimated(121) xor estimated(122) xor estimated(123);
partial_sums(3)(121) <= estimated(632) xor estimated(633) xor estimated(634) xor estimated(635);
partial_sums(3)(122) <= estimated(376) xor estimated(377) xor estimated(378) xor estimated(379);
partial_sums(3)(123) <= estimated(888) xor estimated(889) xor estimated(890) xor estimated(891);
partial_sums(3)(124) <= estimated(248) xor estimated(249) xor estimated(250) xor estimated(251);
partial_sums(3)(125) <= estimated(760) xor estimated(761) xor estimated(762) xor estimated(763);
partial_sums(3)(126) <= estimated(504) xor estimated(505) xor estimated(506) xor estimated(507);
partial_sums(3)(127) <= estimated(1016) xor estimated(1017) xor estimated(1018) xor estimated(1019);
partial_sums(3)(128) <= estimated(2) xor estimated(3);
partial_sums(3)(129) <= estimated(514) xor estimated(515);
partial_sums(3)(130) <= estimated(258) xor estimated(259);
partial_sums(3)(131) <= estimated(770) xor estimated(771);
partial_sums(3)(132) <= estimated(130) xor estimated(131);
partial_sums(3)(133) <= estimated(642) xor estimated(643);
partial_sums(3)(134) <= estimated(386) xor estimated(387);
partial_sums(3)(135) <= estimated(898) xor estimated(899);
partial_sums(3)(136) <= estimated(66) xor estimated(67);
partial_sums(3)(137) <= estimated(578) xor estimated(579);
partial_sums(3)(138) <= estimated(322) xor estimated(323);
partial_sums(3)(139) <= estimated(834) xor estimated(835);
partial_sums(3)(140) <= estimated(194) xor estimated(195);
partial_sums(3)(141) <= estimated(706) xor estimated(707);
partial_sums(3)(142) <= estimated(450) xor estimated(451);
partial_sums(3)(143) <= estimated(962) xor estimated(963);
partial_sums(3)(144) <= estimated(34) xor estimated(35);
partial_sums(3)(145) <= estimated(546) xor estimated(547);
partial_sums(3)(146) <= estimated(290) xor estimated(291);
partial_sums(3)(147) <= estimated(802) xor estimated(803);
partial_sums(3)(148) <= estimated(162) xor estimated(163);
partial_sums(3)(149) <= estimated(674) xor estimated(675);
partial_sums(3)(150) <= estimated(418) xor estimated(419);
partial_sums(3)(151) <= estimated(930) xor estimated(931);
partial_sums(3)(152) <= estimated(98) xor estimated(99);
partial_sums(3)(153) <= estimated(610) xor estimated(611);
partial_sums(3)(154) <= estimated(354) xor estimated(355);
partial_sums(3)(155) <= estimated(866) xor estimated(867);
partial_sums(3)(156) <= estimated(226) xor estimated(227);
partial_sums(3)(157) <= estimated(738) xor estimated(739);
partial_sums(3)(158) <= estimated(482) xor estimated(483);
partial_sums(3)(159) <= estimated(994) xor estimated(995);
partial_sums(3)(160) <= estimated(18) xor estimated(19);
partial_sums(3)(161) <= estimated(530) xor estimated(531);
partial_sums(3)(162) <= estimated(274) xor estimated(275);
partial_sums(3)(163) <= estimated(786) xor estimated(787);
partial_sums(3)(164) <= estimated(146) xor estimated(147);
partial_sums(3)(165) <= estimated(658) xor estimated(659);
partial_sums(3)(166) <= estimated(402) xor estimated(403);
partial_sums(3)(167) <= estimated(914) xor estimated(915);
partial_sums(3)(168) <= estimated(82) xor estimated(83);
partial_sums(3)(169) <= estimated(594) xor estimated(595);
partial_sums(3)(170) <= estimated(338) xor estimated(339);
partial_sums(3)(171) <= estimated(850) xor estimated(851);
partial_sums(3)(172) <= estimated(210) xor estimated(211);
partial_sums(3)(173) <= estimated(722) xor estimated(723);
partial_sums(3)(174) <= estimated(466) xor estimated(467);
partial_sums(3)(175) <= estimated(978) xor estimated(979);
partial_sums(3)(176) <= estimated(50) xor estimated(51);
partial_sums(3)(177) <= estimated(562) xor estimated(563);
partial_sums(3)(178) <= estimated(306) xor estimated(307);
partial_sums(3)(179) <= estimated(818) xor estimated(819);
partial_sums(3)(180) <= estimated(178) xor estimated(179);
partial_sums(3)(181) <= estimated(690) xor estimated(691);
partial_sums(3)(182) <= estimated(434) xor estimated(435);
partial_sums(3)(183) <= estimated(946) xor estimated(947);
partial_sums(3)(184) <= estimated(114) xor estimated(115);
partial_sums(3)(185) <= estimated(626) xor estimated(627);
partial_sums(3)(186) <= estimated(370) xor estimated(371);
partial_sums(3)(187) <= estimated(882) xor estimated(883);
partial_sums(3)(188) <= estimated(242) xor estimated(243);
partial_sums(3)(189) <= estimated(754) xor estimated(755);
partial_sums(3)(190) <= estimated(498) xor estimated(499);
partial_sums(3)(191) <= estimated(1010) xor estimated(1011);
partial_sums(3)(192) <= estimated(10) xor estimated(11);
partial_sums(3)(193) <= estimated(522) xor estimated(523);
partial_sums(3)(194) <= estimated(266) xor estimated(267);
partial_sums(3)(195) <= estimated(778) xor estimated(779);
partial_sums(3)(196) <= estimated(138) xor estimated(139);
partial_sums(3)(197) <= estimated(650) xor estimated(651);
partial_sums(3)(198) <= estimated(394) xor estimated(395);
partial_sums(3)(199) <= estimated(906) xor estimated(907);
partial_sums(3)(200) <= estimated(74) xor estimated(75);
partial_sums(3)(201) <= estimated(586) xor estimated(587);
partial_sums(3)(202) <= estimated(330) xor estimated(331);
partial_sums(3)(203) <= estimated(842) xor estimated(843);
partial_sums(3)(204) <= estimated(202) xor estimated(203);
partial_sums(3)(205) <= estimated(714) xor estimated(715);
partial_sums(3)(206) <= estimated(458) xor estimated(459);
partial_sums(3)(207) <= estimated(970) xor estimated(971);
partial_sums(3)(208) <= estimated(42) xor estimated(43);
partial_sums(3)(209) <= estimated(554) xor estimated(555);
partial_sums(3)(210) <= estimated(298) xor estimated(299);
partial_sums(3)(211) <= estimated(810) xor estimated(811);
partial_sums(3)(212) <= estimated(170) xor estimated(171);
partial_sums(3)(213) <= estimated(682) xor estimated(683);
partial_sums(3)(214) <= estimated(426) xor estimated(427);
partial_sums(3)(215) <= estimated(938) xor estimated(939);
partial_sums(3)(216) <= estimated(106) xor estimated(107);
partial_sums(3)(217) <= estimated(618) xor estimated(619);
partial_sums(3)(218) <= estimated(362) xor estimated(363);
partial_sums(3)(219) <= estimated(874) xor estimated(875);
partial_sums(3)(220) <= estimated(234) xor estimated(235);
partial_sums(3)(221) <= estimated(746) xor estimated(747);
partial_sums(3)(222) <= estimated(490) xor estimated(491);
partial_sums(3)(223) <= estimated(1002) xor estimated(1003);
partial_sums(3)(224) <= estimated(26) xor estimated(27);
partial_sums(3)(225) <= estimated(538) xor estimated(539);
partial_sums(3)(226) <= estimated(282) xor estimated(283);
partial_sums(3)(227) <= estimated(794) xor estimated(795);
partial_sums(3)(228) <= estimated(154) xor estimated(155);
partial_sums(3)(229) <= estimated(666) xor estimated(667);
partial_sums(3)(230) <= estimated(410) xor estimated(411);
partial_sums(3)(231) <= estimated(922) xor estimated(923);
partial_sums(3)(232) <= estimated(90) xor estimated(91);
partial_sums(3)(233) <= estimated(602) xor estimated(603);
partial_sums(3)(234) <= estimated(346) xor estimated(347);
partial_sums(3)(235) <= estimated(858) xor estimated(859);
partial_sums(3)(236) <= estimated(218) xor estimated(219);
partial_sums(3)(237) <= estimated(730) xor estimated(731);
partial_sums(3)(238) <= estimated(474) xor estimated(475);
partial_sums(3)(239) <= estimated(986) xor estimated(987);
partial_sums(3)(240) <= estimated(58) xor estimated(59);
partial_sums(3)(241) <= estimated(570) xor estimated(571);
partial_sums(3)(242) <= estimated(314) xor estimated(315);
partial_sums(3)(243) <= estimated(826) xor estimated(827);
partial_sums(3)(244) <= estimated(186) xor estimated(187);
partial_sums(3)(245) <= estimated(698) xor estimated(699);
partial_sums(3)(246) <= estimated(442) xor estimated(443);
partial_sums(3)(247) <= estimated(954) xor estimated(955);
partial_sums(3)(248) <= estimated(122) xor estimated(123);
partial_sums(3)(249) <= estimated(634) xor estimated(635);
partial_sums(3)(250) <= estimated(378) xor estimated(379);
partial_sums(3)(251) <= estimated(890) xor estimated(891);
partial_sums(3)(252) <= estimated(250) xor estimated(251);
partial_sums(3)(253) <= estimated(762) xor estimated(763);
partial_sums(3)(254) <= estimated(506) xor estimated(507);
partial_sums(3)(255) <= estimated(1018) xor estimated(1019);
partial_sums(3)(256) <= estimated(1) xor estimated(3);
partial_sums(3)(257) <= estimated(513) xor estimated(515);
partial_sums(3)(258) <= estimated(257) xor estimated(259);
partial_sums(3)(259) <= estimated(769) xor estimated(771);
partial_sums(3)(260) <= estimated(129) xor estimated(131);
partial_sums(3)(261) <= estimated(641) xor estimated(643);
partial_sums(3)(262) <= estimated(385) xor estimated(387);
partial_sums(3)(263) <= estimated(897) xor estimated(899);
partial_sums(3)(264) <= estimated(65) xor estimated(67);
partial_sums(3)(265) <= estimated(577) xor estimated(579);
partial_sums(3)(266) <= estimated(321) xor estimated(323);
partial_sums(3)(267) <= estimated(833) xor estimated(835);
partial_sums(3)(268) <= estimated(193) xor estimated(195);
partial_sums(3)(269) <= estimated(705) xor estimated(707);
partial_sums(3)(270) <= estimated(449) xor estimated(451);
partial_sums(3)(271) <= estimated(961) xor estimated(963);
partial_sums(3)(272) <= estimated(33) xor estimated(35);
partial_sums(3)(273) <= estimated(545) xor estimated(547);
partial_sums(3)(274) <= estimated(289) xor estimated(291);
partial_sums(3)(275) <= estimated(801) xor estimated(803);
partial_sums(3)(276) <= estimated(161) xor estimated(163);
partial_sums(3)(277) <= estimated(673) xor estimated(675);
partial_sums(3)(278) <= estimated(417) xor estimated(419);
partial_sums(3)(279) <= estimated(929) xor estimated(931);
partial_sums(3)(280) <= estimated(97) xor estimated(99);
partial_sums(3)(281) <= estimated(609) xor estimated(611);
partial_sums(3)(282) <= estimated(353) xor estimated(355);
partial_sums(3)(283) <= estimated(865) xor estimated(867);
partial_sums(3)(284) <= estimated(225) xor estimated(227);
partial_sums(3)(285) <= estimated(737) xor estimated(739);
partial_sums(3)(286) <= estimated(481) xor estimated(483);
partial_sums(3)(287) <= estimated(993) xor estimated(995);
partial_sums(3)(288) <= estimated(17) xor estimated(19);
partial_sums(3)(289) <= estimated(529) xor estimated(531);
partial_sums(3)(290) <= estimated(273) xor estimated(275);
partial_sums(3)(291) <= estimated(785) xor estimated(787);
partial_sums(3)(292) <= estimated(145) xor estimated(147);
partial_sums(3)(293) <= estimated(657) xor estimated(659);
partial_sums(3)(294) <= estimated(401) xor estimated(403);
partial_sums(3)(295) <= estimated(913) xor estimated(915);
partial_sums(3)(296) <= estimated(81) xor estimated(83);
partial_sums(3)(297) <= estimated(593) xor estimated(595);
partial_sums(3)(298) <= estimated(337) xor estimated(339);
partial_sums(3)(299) <= estimated(849) xor estimated(851);
partial_sums(3)(300) <= estimated(209) xor estimated(211);
partial_sums(3)(301) <= estimated(721) xor estimated(723);
partial_sums(3)(302) <= estimated(465) xor estimated(467);
partial_sums(3)(303) <= estimated(977) xor estimated(979);
partial_sums(3)(304) <= estimated(49) xor estimated(51);
partial_sums(3)(305) <= estimated(561) xor estimated(563);
partial_sums(3)(306) <= estimated(305) xor estimated(307);
partial_sums(3)(307) <= estimated(817) xor estimated(819);
partial_sums(3)(308) <= estimated(177) xor estimated(179);
partial_sums(3)(309) <= estimated(689) xor estimated(691);
partial_sums(3)(310) <= estimated(433) xor estimated(435);
partial_sums(3)(311) <= estimated(945) xor estimated(947);
partial_sums(3)(312) <= estimated(113) xor estimated(115);
partial_sums(3)(313) <= estimated(625) xor estimated(627);
partial_sums(3)(314) <= estimated(369) xor estimated(371);
partial_sums(3)(315) <= estimated(881) xor estimated(883);
partial_sums(3)(316) <= estimated(241) xor estimated(243);
partial_sums(3)(317) <= estimated(753) xor estimated(755);
partial_sums(3)(318) <= estimated(497) xor estimated(499);
partial_sums(3)(319) <= estimated(1009) xor estimated(1011);
partial_sums(3)(320) <= estimated(9) xor estimated(11);
partial_sums(3)(321) <= estimated(521) xor estimated(523);
partial_sums(3)(322) <= estimated(265) xor estimated(267);
partial_sums(3)(323) <= estimated(777) xor estimated(779);
partial_sums(3)(324) <= estimated(137) xor estimated(139);
partial_sums(3)(325) <= estimated(649) xor estimated(651);
partial_sums(3)(326) <= estimated(393) xor estimated(395);
partial_sums(3)(327) <= estimated(905) xor estimated(907);
partial_sums(3)(328) <= estimated(73) xor estimated(75);
partial_sums(3)(329) <= estimated(585) xor estimated(587);
partial_sums(3)(330) <= estimated(329) xor estimated(331);
partial_sums(3)(331) <= estimated(841) xor estimated(843);
partial_sums(3)(332) <= estimated(201) xor estimated(203);
partial_sums(3)(333) <= estimated(713) xor estimated(715);
partial_sums(3)(334) <= estimated(457) xor estimated(459);
partial_sums(3)(335) <= estimated(969) xor estimated(971);
partial_sums(3)(336) <= estimated(41) xor estimated(43);
partial_sums(3)(337) <= estimated(553) xor estimated(555);
partial_sums(3)(338) <= estimated(297) xor estimated(299);
partial_sums(3)(339) <= estimated(809) xor estimated(811);
partial_sums(3)(340) <= estimated(169) xor estimated(171);
partial_sums(3)(341) <= estimated(681) xor estimated(683);
partial_sums(3)(342) <= estimated(425) xor estimated(427);
partial_sums(3)(343) <= estimated(937) xor estimated(939);
partial_sums(3)(344) <= estimated(105) xor estimated(107);
partial_sums(3)(345) <= estimated(617) xor estimated(619);
partial_sums(3)(346) <= estimated(361) xor estimated(363);
partial_sums(3)(347) <= estimated(873) xor estimated(875);
partial_sums(3)(348) <= estimated(233) xor estimated(235);
partial_sums(3)(349) <= estimated(745) xor estimated(747);
partial_sums(3)(350) <= estimated(489) xor estimated(491);
partial_sums(3)(351) <= estimated(1001) xor estimated(1003);
partial_sums(3)(352) <= estimated(25) xor estimated(27);
partial_sums(3)(353) <= estimated(537) xor estimated(539);
partial_sums(3)(354) <= estimated(281) xor estimated(283);
partial_sums(3)(355) <= estimated(793) xor estimated(795);
partial_sums(3)(356) <= estimated(153) xor estimated(155);
partial_sums(3)(357) <= estimated(665) xor estimated(667);
partial_sums(3)(358) <= estimated(409) xor estimated(411);
partial_sums(3)(359) <= estimated(921) xor estimated(923);
partial_sums(3)(360) <= estimated(89) xor estimated(91);
partial_sums(3)(361) <= estimated(601) xor estimated(603);
partial_sums(3)(362) <= estimated(345) xor estimated(347);
partial_sums(3)(363) <= estimated(857) xor estimated(859);
partial_sums(3)(364) <= estimated(217) xor estimated(219);
partial_sums(3)(365) <= estimated(729) xor estimated(731);
partial_sums(3)(366) <= estimated(473) xor estimated(475);
partial_sums(3)(367) <= estimated(985) xor estimated(987);
partial_sums(3)(368) <= estimated(57) xor estimated(59);
partial_sums(3)(369) <= estimated(569) xor estimated(571);
partial_sums(3)(370) <= estimated(313) xor estimated(315);
partial_sums(3)(371) <= estimated(825) xor estimated(827);
partial_sums(3)(372) <= estimated(185) xor estimated(187);
partial_sums(3)(373) <= estimated(697) xor estimated(699);
partial_sums(3)(374) <= estimated(441) xor estimated(443);
partial_sums(3)(375) <= estimated(953) xor estimated(955);
partial_sums(3)(376) <= estimated(121) xor estimated(123);
partial_sums(3)(377) <= estimated(633) xor estimated(635);
partial_sums(3)(378) <= estimated(377) xor estimated(379);
partial_sums(3)(379) <= estimated(889) xor estimated(891);
partial_sums(3)(380) <= estimated(249) xor estimated(251);
partial_sums(3)(381) <= estimated(761) xor estimated(763);
partial_sums(3)(382) <= estimated(505) xor estimated(507);
partial_sums(3)(383) <= estimated(1017) xor estimated(1019);
partial_sums(3)(384) <= estimated(3);
partial_sums(3)(385) <= estimated(515);
partial_sums(3)(386) <= estimated(259);
partial_sums(3)(387) <= estimated(771);
partial_sums(3)(388) <= estimated(131);
partial_sums(3)(389) <= estimated(643);
partial_sums(3)(390) <= estimated(387);
partial_sums(3)(391) <= estimated(899);
partial_sums(3)(392) <= estimated(67);
partial_sums(3)(393) <= estimated(579);
partial_sums(3)(394) <= estimated(323);
partial_sums(3)(395) <= estimated(835);
partial_sums(3)(396) <= estimated(195);
partial_sums(3)(397) <= estimated(707);
partial_sums(3)(398) <= estimated(451);
partial_sums(3)(399) <= estimated(963);
partial_sums(3)(400) <= estimated(35);
partial_sums(3)(401) <= estimated(547);
partial_sums(3)(402) <= estimated(291);
partial_sums(3)(403) <= estimated(803);
partial_sums(3)(404) <= estimated(163);
partial_sums(3)(405) <= estimated(675);
partial_sums(3)(406) <= estimated(419);
partial_sums(3)(407) <= estimated(931);
partial_sums(3)(408) <= estimated(99);
partial_sums(3)(409) <= estimated(611);
partial_sums(3)(410) <= estimated(355);
partial_sums(3)(411) <= estimated(867);
partial_sums(3)(412) <= estimated(227);
partial_sums(3)(413) <= estimated(739);
partial_sums(3)(414) <= estimated(483);
partial_sums(3)(415) <= estimated(995);
partial_sums(3)(416) <= estimated(19);
partial_sums(3)(417) <= estimated(531);
partial_sums(3)(418) <= estimated(275);
partial_sums(3)(419) <= estimated(787);
partial_sums(3)(420) <= estimated(147);
partial_sums(3)(421) <= estimated(659);
partial_sums(3)(422) <= estimated(403);
partial_sums(3)(423) <= estimated(915);
partial_sums(3)(424) <= estimated(83);
partial_sums(3)(425) <= estimated(595);
partial_sums(3)(426) <= estimated(339);
partial_sums(3)(427) <= estimated(851);
partial_sums(3)(428) <= estimated(211);
partial_sums(3)(429) <= estimated(723);
partial_sums(3)(430) <= estimated(467);
partial_sums(3)(431) <= estimated(979);
partial_sums(3)(432) <= estimated(51);
partial_sums(3)(433) <= estimated(563);
partial_sums(3)(434) <= estimated(307);
partial_sums(3)(435) <= estimated(819);
partial_sums(3)(436) <= estimated(179);
partial_sums(3)(437) <= estimated(691);
partial_sums(3)(438) <= estimated(435);
partial_sums(3)(439) <= estimated(947);
partial_sums(3)(440) <= estimated(115);
partial_sums(3)(441) <= estimated(627);
partial_sums(3)(442) <= estimated(371);
partial_sums(3)(443) <= estimated(883);
partial_sums(3)(444) <= estimated(243);
partial_sums(3)(445) <= estimated(755);
partial_sums(3)(446) <= estimated(499);
partial_sums(3)(447) <= estimated(1011);
partial_sums(3)(448) <= estimated(11);
partial_sums(3)(449) <= estimated(523);
partial_sums(3)(450) <= estimated(267);
partial_sums(3)(451) <= estimated(779);
partial_sums(3)(452) <= estimated(139);
partial_sums(3)(453) <= estimated(651);
partial_sums(3)(454) <= estimated(395);
partial_sums(3)(455) <= estimated(907);
partial_sums(3)(456) <= estimated(75);
partial_sums(3)(457) <= estimated(587);
partial_sums(3)(458) <= estimated(331);
partial_sums(3)(459) <= estimated(843);
partial_sums(3)(460) <= estimated(203);
partial_sums(3)(461) <= estimated(715);
partial_sums(3)(462) <= estimated(459);
partial_sums(3)(463) <= estimated(971);
partial_sums(3)(464) <= estimated(43);
partial_sums(3)(465) <= estimated(555);
partial_sums(3)(466) <= estimated(299);
partial_sums(3)(467) <= estimated(811);
partial_sums(3)(468) <= estimated(171);
partial_sums(3)(469) <= estimated(683);
partial_sums(3)(470) <= estimated(427);
partial_sums(3)(471) <= estimated(939);
partial_sums(3)(472) <= estimated(107);
partial_sums(3)(473) <= estimated(619);
partial_sums(3)(474) <= estimated(363);
partial_sums(3)(475) <= estimated(875);
partial_sums(3)(476) <= estimated(235);
partial_sums(3)(477) <= estimated(747);
partial_sums(3)(478) <= estimated(491);
partial_sums(3)(479) <= estimated(1003);
partial_sums(3)(480) <= estimated(27);
partial_sums(3)(481) <= estimated(539);
partial_sums(3)(482) <= estimated(283);
partial_sums(3)(483) <= estimated(795);
partial_sums(3)(484) <= estimated(155);
partial_sums(3)(485) <= estimated(667);
partial_sums(3)(486) <= estimated(411);
partial_sums(3)(487) <= estimated(923);
partial_sums(3)(488) <= estimated(91);
partial_sums(3)(489) <= estimated(603);
partial_sums(3)(490) <= estimated(347);
partial_sums(3)(491) <= estimated(859);
partial_sums(3)(492) <= estimated(219);
partial_sums(3)(493) <= estimated(731);
partial_sums(3)(494) <= estimated(475);
partial_sums(3)(495) <= estimated(987);
partial_sums(3)(496) <= estimated(59);
partial_sums(3)(497) <= estimated(571);
partial_sums(3)(498) <= estimated(315);
partial_sums(3)(499) <= estimated(827);
partial_sums(3)(500) <= estimated(187);
partial_sums(3)(501) <= estimated(699);
partial_sums(3)(502) <= estimated(443);
partial_sums(3)(503) <= estimated(955);
partial_sums(3)(504) <= estimated(123);
partial_sums(3)(505) <= estimated(635);
partial_sums(3)(506) <= estimated(379);
partial_sums(3)(507) <= estimated(891);
partial_sums(3)(508) <= estimated(251);
partial_sums(3)(509) <= estimated(763);
partial_sums(3)(510) <= estimated(507);
partial_sums(3)(511) <= estimated(1019);
partial_sums(4)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7);
partial_sums(4)(1) <= estimated(512) xor estimated(513) xor estimated(514) xor estimated(515) xor estimated(516) xor estimated(517) xor estimated(518) xor estimated(519);
partial_sums(4)(2) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263);
partial_sums(4)(3) <= estimated(768) xor estimated(769) xor estimated(770) xor estimated(771) xor estimated(772) xor estimated(773) xor estimated(774) xor estimated(775);
partial_sums(4)(4) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135);
partial_sums(4)(5) <= estimated(640) xor estimated(641) xor estimated(642) xor estimated(643) xor estimated(644) xor estimated(645) xor estimated(646) xor estimated(647);
partial_sums(4)(6) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391);
partial_sums(4)(7) <= estimated(896) xor estimated(897) xor estimated(898) xor estimated(899) xor estimated(900) xor estimated(901) xor estimated(902) xor estimated(903);
partial_sums(4)(8) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71);
partial_sums(4)(9) <= estimated(576) xor estimated(577) xor estimated(578) xor estimated(579) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583);
partial_sums(4)(10) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327);
partial_sums(4)(11) <= estimated(832) xor estimated(833) xor estimated(834) xor estimated(835) xor estimated(836) xor estimated(837) xor estimated(838) xor estimated(839);
partial_sums(4)(12) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199);
partial_sums(4)(13) <= estimated(704) xor estimated(705) xor estimated(706) xor estimated(707) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711);
partial_sums(4)(14) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455);
partial_sums(4)(15) <= estimated(960) xor estimated(961) xor estimated(962) xor estimated(963) xor estimated(964) xor estimated(965) xor estimated(966) xor estimated(967);
partial_sums(4)(16) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39);
partial_sums(4)(17) <= estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551);
partial_sums(4)(18) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295);
partial_sums(4)(19) <= estimated(800) xor estimated(801) xor estimated(802) xor estimated(803) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807);
partial_sums(4)(20) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167);
partial_sums(4)(21) <= estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679);
partial_sums(4)(22) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423);
partial_sums(4)(23) <= estimated(928) xor estimated(929) xor estimated(930) xor estimated(931) xor estimated(932) xor estimated(933) xor estimated(934) xor estimated(935);
partial_sums(4)(24) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103);
partial_sums(4)(25) <= estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615);
partial_sums(4)(26) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359);
partial_sums(4)(27) <= estimated(864) xor estimated(865) xor estimated(866) xor estimated(867) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871);
partial_sums(4)(28) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231);
partial_sums(4)(29) <= estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743);
partial_sums(4)(30) <= estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487);
partial_sums(4)(31) <= estimated(992) xor estimated(993) xor estimated(994) xor estimated(995) xor estimated(996) xor estimated(997) xor estimated(998) xor estimated(999);
partial_sums(4)(32) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23);
partial_sums(4)(33) <= estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535);
partial_sums(4)(34) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279);
partial_sums(4)(35) <= estimated(784) xor estimated(785) xor estimated(786) xor estimated(787) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791);
partial_sums(4)(36) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151);
partial_sums(4)(37) <= estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663);
partial_sums(4)(38) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407);
partial_sums(4)(39) <= estimated(912) xor estimated(913) xor estimated(914) xor estimated(915) xor estimated(916) xor estimated(917) xor estimated(918) xor estimated(919);
partial_sums(4)(40) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87);
partial_sums(4)(41) <= estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599);
partial_sums(4)(42) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343);
partial_sums(4)(43) <= estimated(848) xor estimated(849) xor estimated(850) xor estimated(851) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855);
partial_sums(4)(44) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215);
partial_sums(4)(45) <= estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727);
partial_sums(4)(46) <= estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471);
partial_sums(4)(47) <= estimated(976) xor estimated(977) xor estimated(978) xor estimated(979) xor estimated(980) xor estimated(981) xor estimated(982) xor estimated(983);
partial_sums(4)(48) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55);
partial_sums(4)(49) <= estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567);
partial_sums(4)(50) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311);
partial_sums(4)(51) <= estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823);
partial_sums(4)(52) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183);
partial_sums(4)(53) <= estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695);
partial_sums(4)(54) <= estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439);
partial_sums(4)(55) <= estimated(944) xor estimated(945) xor estimated(946) xor estimated(947) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951);
partial_sums(4)(56) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119);
partial_sums(4)(57) <= estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631);
partial_sums(4)(58) <= estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375);
partial_sums(4)(59) <= estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887);
partial_sums(4)(60) <= estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247);
partial_sums(4)(61) <= estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759);
partial_sums(4)(62) <= estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503);
partial_sums(4)(63) <= estimated(1008) xor estimated(1009) xor estimated(1010) xor estimated(1011) xor estimated(1012) xor estimated(1013) xor estimated(1014) xor estimated(1015);
partial_sums(4)(64) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7);
partial_sums(4)(65) <= estimated(516) xor estimated(517) xor estimated(518) xor estimated(519);
partial_sums(4)(66) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263);
partial_sums(4)(67) <= estimated(772) xor estimated(773) xor estimated(774) xor estimated(775);
partial_sums(4)(68) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135);
partial_sums(4)(69) <= estimated(644) xor estimated(645) xor estimated(646) xor estimated(647);
partial_sums(4)(70) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391);
partial_sums(4)(71) <= estimated(900) xor estimated(901) xor estimated(902) xor estimated(903);
partial_sums(4)(72) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71);
partial_sums(4)(73) <= estimated(580) xor estimated(581) xor estimated(582) xor estimated(583);
partial_sums(4)(74) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327);
partial_sums(4)(75) <= estimated(836) xor estimated(837) xor estimated(838) xor estimated(839);
partial_sums(4)(76) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199);
partial_sums(4)(77) <= estimated(708) xor estimated(709) xor estimated(710) xor estimated(711);
partial_sums(4)(78) <= estimated(452) xor estimated(453) xor estimated(454) xor estimated(455);
partial_sums(4)(79) <= estimated(964) xor estimated(965) xor estimated(966) xor estimated(967);
partial_sums(4)(80) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39);
partial_sums(4)(81) <= estimated(548) xor estimated(549) xor estimated(550) xor estimated(551);
partial_sums(4)(82) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295);
partial_sums(4)(83) <= estimated(804) xor estimated(805) xor estimated(806) xor estimated(807);
partial_sums(4)(84) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167);
partial_sums(4)(85) <= estimated(676) xor estimated(677) xor estimated(678) xor estimated(679);
partial_sums(4)(86) <= estimated(420) xor estimated(421) xor estimated(422) xor estimated(423);
partial_sums(4)(87) <= estimated(932) xor estimated(933) xor estimated(934) xor estimated(935);
partial_sums(4)(88) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103);
partial_sums(4)(89) <= estimated(612) xor estimated(613) xor estimated(614) xor estimated(615);
partial_sums(4)(90) <= estimated(356) xor estimated(357) xor estimated(358) xor estimated(359);
partial_sums(4)(91) <= estimated(868) xor estimated(869) xor estimated(870) xor estimated(871);
partial_sums(4)(92) <= estimated(228) xor estimated(229) xor estimated(230) xor estimated(231);
partial_sums(4)(93) <= estimated(740) xor estimated(741) xor estimated(742) xor estimated(743);
partial_sums(4)(94) <= estimated(484) xor estimated(485) xor estimated(486) xor estimated(487);
partial_sums(4)(95) <= estimated(996) xor estimated(997) xor estimated(998) xor estimated(999);
partial_sums(4)(96) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23);
partial_sums(4)(97) <= estimated(532) xor estimated(533) xor estimated(534) xor estimated(535);
partial_sums(4)(98) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279);
partial_sums(4)(99) <= estimated(788) xor estimated(789) xor estimated(790) xor estimated(791);
partial_sums(4)(100) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151);
partial_sums(4)(101) <= estimated(660) xor estimated(661) xor estimated(662) xor estimated(663);
partial_sums(4)(102) <= estimated(404) xor estimated(405) xor estimated(406) xor estimated(407);
partial_sums(4)(103) <= estimated(916) xor estimated(917) xor estimated(918) xor estimated(919);
partial_sums(4)(104) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87);
partial_sums(4)(105) <= estimated(596) xor estimated(597) xor estimated(598) xor estimated(599);
partial_sums(4)(106) <= estimated(340) xor estimated(341) xor estimated(342) xor estimated(343);
partial_sums(4)(107) <= estimated(852) xor estimated(853) xor estimated(854) xor estimated(855);
partial_sums(4)(108) <= estimated(212) xor estimated(213) xor estimated(214) xor estimated(215);
partial_sums(4)(109) <= estimated(724) xor estimated(725) xor estimated(726) xor estimated(727);
partial_sums(4)(110) <= estimated(468) xor estimated(469) xor estimated(470) xor estimated(471);
partial_sums(4)(111) <= estimated(980) xor estimated(981) xor estimated(982) xor estimated(983);
partial_sums(4)(112) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55);
partial_sums(4)(113) <= estimated(564) xor estimated(565) xor estimated(566) xor estimated(567);
partial_sums(4)(114) <= estimated(308) xor estimated(309) xor estimated(310) xor estimated(311);
partial_sums(4)(115) <= estimated(820) xor estimated(821) xor estimated(822) xor estimated(823);
partial_sums(4)(116) <= estimated(180) xor estimated(181) xor estimated(182) xor estimated(183);
partial_sums(4)(117) <= estimated(692) xor estimated(693) xor estimated(694) xor estimated(695);
partial_sums(4)(118) <= estimated(436) xor estimated(437) xor estimated(438) xor estimated(439);
partial_sums(4)(119) <= estimated(948) xor estimated(949) xor estimated(950) xor estimated(951);
partial_sums(4)(120) <= estimated(116) xor estimated(117) xor estimated(118) xor estimated(119);
partial_sums(4)(121) <= estimated(628) xor estimated(629) xor estimated(630) xor estimated(631);
partial_sums(4)(122) <= estimated(372) xor estimated(373) xor estimated(374) xor estimated(375);
partial_sums(4)(123) <= estimated(884) xor estimated(885) xor estimated(886) xor estimated(887);
partial_sums(4)(124) <= estimated(244) xor estimated(245) xor estimated(246) xor estimated(247);
partial_sums(4)(125) <= estimated(756) xor estimated(757) xor estimated(758) xor estimated(759);
partial_sums(4)(126) <= estimated(500) xor estimated(501) xor estimated(502) xor estimated(503);
partial_sums(4)(127) <= estimated(1012) xor estimated(1013) xor estimated(1014) xor estimated(1015);
partial_sums(4)(128) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7);
partial_sums(4)(129) <= estimated(514) xor estimated(515) xor estimated(518) xor estimated(519);
partial_sums(4)(130) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263);
partial_sums(4)(131) <= estimated(770) xor estimated(771) xor estimated(774) xor estimated(775);
partial_sums(4)(132) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135);
partial_sums(4)(133) <= estimated(642) xor estimated(643) xor estimated(646) xor estimated(647);
partial_sums(4)(134) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391);
partial_sums(4)(135) <= estimated(898) xor estimated(899) xor estimated(902) xor estimated(903);
partial_sums(4)(136) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71);
partial_sums(4)(137) <= estimated(578) xor estimated(579) xor estimated(582) xor estimated(583);
partial_sums(4)(138) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327);
partial_sums(4)(139) <= estimated(834) xor estimated(835) xor estimated(838) xor estimated(839);
partial_sums(4)(140) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199);
partial_sums(4)(141) <= estimated(706) xor estimated(707) xor estimated(710) xor estimated(711);
partial_sums(4)(142) <= estimated(450) xor estimated(451) xor estimated(454) xor estimated(455);
partial_sums(4)(143) <= estimated(962) xor estimated(963) xor estimated(966) xor estimated(967);
partial_sums(4)(144) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39);
partial_sums(4)(145) <= estimated(546) xor estimated(547) xor estimated(550) xor estimated(551);
partial_sums(4)(146) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295);
partial_sums(4)(147) <= estimated(802) xor estimated(803) xor estimated(806) xor estimated(807);
partial_sums(4)(148) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167);
partial_sums(4)(149) <= estimated(674) xor estimated(675) xor estimated(678) xor estimated(679);
partial_sums(4)(150) <= estimated(418) xor estimated(419) xor estimated(422) xor estimated(423);
partial_sums(4)(151) <= estimated(930) xor estimated(931) xor estimated(934) xor estimated(935);
partial_sums(4)(152) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103);
partial_sums(4)(153) <= estimated(610) xor estimated(611) xor estimated(614) xor estimated(615);
partial_sums(4)(154) <= estimated(354) xor estimated(355) xor estimated(358) xor estimated(359);
partial_sums(4)(155) <= estimated(866) xor estimated(867) xor estimated(870) xor estimated(871);
partial_sums(4)(156) <= estimated(226) xor estimated(227) xor estimated(230) xor estimated(231);
partial_sums(4)(157) <= estimated(738) xor estimated(739) xor estimated(742) xor estimated(743);
partial_sums(4)(158) <= estimated(482) xor estimated(483) xor estimated(486) xor estimated(487);
partial_sums(4)(159) <= estimated(994) xor estimated(995) xor estimated(998) xor estimated(999);
partial_sums(4)(160) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23);
partial_sums(4)(161) <= estimated(530) xor estimated(531) xor estimated(534) xor estimated(535);
partial_sums(4)(162) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279);
partial_sums(4)(163) <= estimated(786) xor estimated(787) xor estimated(790) xor estimated(791);
partial_sums(4)(164) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151);
partial_sums(4)(165) <= estimated(658) xor estimated(659) xor estimated(662) xor estimated(663);
partial_sums(4)(166) <= estimated(402) xor estimated(403) xor estimated(406) xor estimated(407);
partial_sums(4)(167) <= estimated(914) xor estimated(915) xor estimated(918) xor estimated(919);
partial_sums(4)(168) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87);
partial_sums(4)(169) <= estimated(594) xor estimated(595) xor estimated(598) xor estimated(599);
partial_sums(4)(170) <= estimated(338) xor estimated(339) xor estimated(342) xor estimated(343);
partial_sums(4)(171) <= estimated(850) xor estimated(851) xor estimated(854) xor estimated(855);
partial_sums(4)(172) <= estimated(210) xor estimated(211) xor estimated(214) xor estimated(215);
partial_sums(4)(173) <= estimated(722) xor estimated(723) xor estimated(726) xor estimated(727);
partial_sums(4)(174) <= estimated(466) xor estimated(467) xor estimated(470) xor estimated(471);
partial_sums(4)(175) <= estimated(978) xor estimated(979) xor estimated(982) xor estimated(983);
partial_sums(4)(176) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55);
partial_sums(4)(177) <= estimated(562) xor estimated(563) xor estimated(566) xor estimated(567);
partial_sums(4)(178) <= estimated(306) xor estimated(307) xor estimated(310) xor estimated(311);
partial_sums(4)(179) <= estimated(818) xor estimated(819) xor estimated(822) xor estimated(823);
partial_sums(4)(180) <= estimated(178) xor estimated(179) xor estimated(182) xor estimated(183);
partial_sums(4)(181) <= estimated(690) xor estimated(691) xor estimated(694) xor estimated(695);
partial_sums(4)(182) <= estimated(434) xor estimated(435) xor estimated(438) xor estimated(439);
partial_sums(4)(183) <= estimated(946) xor estimated(947) xor estimated(950) xor estimated(951);
partial_sums(4)(184) <= estimated(114) xor estimated(115) xor estimated(118) xor estimated(119);
partial_sums(4)(185) <= estimated(626) xor estimated(627) xor estimated(630) xor estimated(631);
partial_sums(4)(186) <= estimated(370) xor estimated(371) xor estimated(374) xor estimated(375);
partial_sums(4)(187) <= estimated(882) xor estimated(883) xor estimated(886) xor estimated(887);
partial_sums(4)(188) <= estimated(242) xor estimated(243) xor estimated(246) xor estimated(247);
partial_sums(4)(189) <= estimated(754) xor estimated(755) xor estimated(758) xor estimated(759);
partial_sums(4)(190) <= estimated(498) xor estimated(499) xor estimated(502) xor estimated(503);
partial_sums(4)(191) <= estimated(1010) xor estimated(1011) xor estimated(1014) xor estimated(1015);
partial_sums(4)(192) <= estimated(6) xor estimated(7);
partial_sums(4)(193) <= estimated(518) xor estimated(519);
partial_sums(4)(194) <= estimated(262) xor estimated(263);
partial_sums(4)(195) <= estimated(774) xor estimated(775);
partial_sums(4)(196) <= estimated(134) xor estimated(135);
partial_sums(4)(197) <= estimated(646) xor estimated(647);
partial_sums(4)(198) <= estimated(390) xor estimated(391);
partial_sums(4)(199) <= estimated(902) xor estimated(903);
partial_sums(4)(200) <= estimated(70) xor estimated(71);
partial_sums(4)(201) <= estimated(582) xor estimated(583);
partial_sums(4)(202) <= estimated(326) xor estimated(327);
partial_sums(4)(203) <= estimated(838) xor estimated(839);
partial_sums(4)(204) <= estimated(198) xor estimated(199);
partial_sums(4)(205) <= estimated(710) xor estimated(711);
partial_sums(4)(206) <= estimated(454) xor estimated(455);
partial_sums(4)(207) <= estimated(966) xor estimated(967);
partial_sums(4)(208) <= estimated(38) xor estimated(39);
partial_sums(4)(209) <= estimated(550) xor estimated(551);
partial_sums(4)(210) <= estimated(294) xor estimated(295);
partial_sums(4)(211) <= estimated(806) xor estimated(807);
partial_sums(4)(212) <= estimated(166) xor estimated(167);
partial_sums(4)(213) <= estimated(678) xor estimated(679);
partial_sums(4)(214) <= estimated(422) xor estimated(423);
partial_sums(4)(215) <= estimated(934) xor estimated(935);
partial_sums(4)(216) <= estimated(102) xor estimated(103);
partial_sums(4)(217) <= estimated(614) xor estimated(615);
partial_sums(4)(218) <= estimated(358) xor estimated(359);
partial_sums(4)(219) <= estimated(870) xor estimated(871);
partial_sums(4)(220) <= estimated(230) xor estimated(231);
partial_sums(4)(221) <= estimated(742) xor estimated(743);
partial_sums(4)(222) <= estimated(486) xor estimated(487);
partial_sums(4)(223) <= estimated(998) xor estimated(999);
partial_sums(4)(224) <= estimated(22) xor estimated(23);
partial_sums(4)(225) <= estimated(534) xor estimated(535);
partial_sums(4)(226) <= estimated(278) xor estimated(279);
partial_sums(4)(227) <= estimated(790) xor estimated(791);
partial_sums(4)(228) <= estimated(150) xor estimated(151);
partial_sums(4)(229) <= estimated(662) xor estimated(663);
partial_sums(4)(230) <= estimated(406) xor estimated(407);
partial_sums(4)(231) <= estimated(918) xor estimated(919);
partial_sums(4)(232) <= estimated(86) xor estimated(87);
partial_sums(4)(233) <= estimated(598) xor estimated(599);
partial_sums(4)(234) <= estimated(342) xor estimated(343);
partial_sums(4)(235) <= estimated(854) xor estimated(855);
partial_sums(4)(236) <= estimated(214) xor estimated(215);
partial_sums(4)(237) <= estimated(726) xor estimated(727);
partial_sums(4)(238) <= estimated(470) xor estimated(471);
partial_sums(4)(239) <= estimated(982) xor estimated(983);
partial_sums(4)(240) <= estimated(54) xor estimated(55);
partial_sums(4)(241) <= estimated(566) xor estimated(567);
partial_sums(4)(242) <= estimated(310) xor estimated(311);
partial_sums(4)(243) <= estimated(822) xor estimated(823);
partial_sums(4)(244) <= estimated(182) xor estimated(183);
partial_sums(4)(245) <= estimated(694) xor estimated(695);
partial_sums(4)(246) <= estimated(438) xor estimated(439);
partial_sums(4)(247) <= estimated(950) xor estimated(951);
partial_sums(4)(248) <= estimated(118) xor estimated(119);
partial_sums(4)(249) <= estimated(630) xor estimated(631);
partial_sums(4)(250) <= estimated(374) xor estimated(375);
partial_sums(4)(251) <= estimated(886) xor estimated(887);
partial_sums(4)(252) <= estimated(246) xor estimated(247);
partial_sums(4)(253) <= estimated(758) xor estimated(759);
partial_sums(4)(254) <= estimated(502) xor estimated(503);
partial_sums(4)(255) <= estimated(1014) xor estimated(1015);
partial_sums(4)(256) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7);
partial_sums(4)(257) <= estimated(513) xor estimated(515) xor estimated(517) xor estimated(519);
partial_sums(4)(258) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263);
partial_sums(4)(259) <= estimated(769) xor estimated(771) xor estimated(773) xor estimated(775);
partial_sums(4)(260) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135);
partial_sums(4)(261) <= estimated(641) xor estimated(643) xor estimated(645) xor estimated(647);
partial_sums(4)(262) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391);
partial_sums(4)(263) <= estimated(897) xor estimated(899) xor estimated(901) xor estimated(903);
partial_sums(4)(264) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71);
partial_sums(4)(265) <= estimated(577) xor estimated(579) xor estimated(581) xor estimated(583);
partial_sums(4)(266) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327);
partial_sums(4)(267) <= estimated(833) xor estimated(835) xor estimated(837) xor estimated(839);
partial_sums(4)(268) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199);
partial_sums(4)(269) <= estimated(705) xor estimated(707) xor estimated(709) xor estimated(711);
partial_sums(4)(270) <= estimated(449) xor estimated(451) xor estimated(453) xor estimated(455);
partial_sums(4)(271) <= estimated(961) xor estimated(963) xor estimated(965) xor estimated(967);
partial_sums(4)(272) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39);
partial_sums(4)(273) <= estimated(545) xor estimated(547) xor estimated(549) xor estimated(551);
partial_sums(4)(274) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295);
partial_sums(4)(275) <= estimated(801) xor estimated(803) xor estimated(805) xor estimated(807);
partial_sums(4)(276) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167);
partial_sums(4)(277) <= estimated(673) xor estimated(675) xor estimated(677) xor estimated(679);
partial_sums(4)(278) <= estimated(417) xor estimated(419) xor estimated(421) xor estimated(423);
partial_sums(4)(279) <= estimated(929) xor estimated(931) xor estimated(933) xor estimated(935);
partial_sums(4)(280) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103);
partial_sums(4)(281) <= estimated(609) xor estimated(611) xor estimated(613) xor estimated(615);
partial_sums(4)(282) <= estimated(353) xor estimated(355) xor estimated(357) xor estimated(359);
partial_sums(4)(283) <= estimated(865) xor estimated(867) xor estimated(869) xor estimated(871);
partial_sums(4)(284) <= estimated(225) xor estimated(227) xor estimated(229) xor estimated(231);
partial_sums(4)(285) <= estimated(737) xor estimated(739) xor estimated(741) xor estimated(743);
partial_sums(4)(286) <= estimated(481) xor estimated(483) xor estimated(485) xor estimated(487);
partial_sums(4)(287) <= estimated(993) xor estimated(995) xor estimated(997) xor estimated(999);
partial_sums(4)(288) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23);
partial_sums(4)(289) <= estimated(529) xor estimated(531) xor estimated(533) xor estimated(535);
partial_sums(4)(290) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279);
partial_sums(4)(291) <= estimated(785) xor estimated(787) xor estimated(789) xor estimated(791);
partial_sums(4)(292) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151);
partial_sums(4)(293) <= estimated(657) xor estimated(659) xor estimated(661) xor estimated(663);
partial_sums(4)(294) <= estimated(401) xor estimated(403) xor estimated(405) xor estimated(407);
partial_sums(4)(295) <= estimated(913) xor estimated(915) xor estimated(917) xor estimated(919);
partial_sums(4)(296) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87);
partial_sums(4)(297) <= estimated(593) xor estimated(595) xor estimated(597) xor estimated(599);
partial_sums(4)(298) <= estimated(337) xor estimated(339) xor estimated(341) xor estimated(343);
partial_sums(4)(299) <= estimated(849) xor estimated(851) xor estimated(853) xor estimated(855);
partial_sums(4)(300) <= estimated(209) xor estimated(211) xor estimated(213) xor estimated(215);
partial_sums(4)(301) <= estimated(721) xor estimated(723) xor estimated(725) xor estimated(727);
partial_sums(4)(302) <= estimated(465) xor estimated(467) xor estimated(469) xor estimated(471);
partial_sums(4)(303) <= estimated(977) xor estimated(979) xor estimated(981) xor estimated(983);
partial_sums(4)(304) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55);
partial_sums(4)(305) <= estimated(561) xor estimated(563) xor estimated(565) xor estimated(567);
partial_sums(4)(306) <= estimated(305) xor estimated(307) xor estimated(309) xor estimated(311);
partial_sums(4)(307) <= estimated(817) xor estimated(819) xor estimated(821) xor estimated(823);
partial_sums(4)(308) <= estimated(177) xor estimated(179) xor estimated(181) xor estimated(183);
partial_sums(4)(309) <= estimated(689) xor estimated(691) xor estimated(693) xor estimated(695);
partial_sums(4)(310) <= estimated(433) xor estimated(435) xor estimated(437) xor estimated(439);
partial_sums(4)(311) <= estimated(945) xor estimated(947) xor estimated(949) xor estimated(951);
partial_sums(4)(312) <= estimated(113) xor estimated(115) xor estimated(117) xor estimated(119);
partial_sums(4)(313) <= estimated(625) xor estimated(627) xor estimated(629) xor estimated(631);
partial_sums(4)(314) <= estimated(369) xor estimated(371) xor estimated(373) xor estimated(375);
partial_sums(4)(315) <= estimated(881) xor estimated(883) xor estimated(885) xor estimated(887);
partial_sums(4)(316) <= estimated(241) xor estimated(243) xor estimated(245) xor estimated(247);
partial_sums(4)(317) <= estimated(753) xor estimated(755) xor estimated(757) xor estimated(759);
partial_sums(4)(318) <= estimated(497) xor estimated(499) xor estimated(501) xor estimated(503);
partial_sums(4)(319) <= estimated(1009) xor estimated(1011) xor estimated(1013) xor estimated(1015);
partial_sums(4)(320) <= estimated(5) xor estimated(7);
partial_sums(4)(321) <= estimated(517) xor estimated(519);
partial_sums(4)(322) <= estimated(261) xor estimated(263);
partial_sums(4)(323) <= estimated(773) xor estimated(775);
partial_sums(4)(324) <= estimated(133) xor estimated(135);
partial_sums(4)(325) <= estimated(645) xor estimated(647);
partial_sums(4)(326) <= estimated(389) xor estimated(391);
partial_sums(4)(327) <= estimated(901) xor estimated(903);
partial_sums(4)(328) <= estimated(69) xor estimated(71);
partial_sums(4)(329) <= estimated(581) xor estimated(583);
partial_sums(4)(330) <= estimated(325) xor estimated(327);
partial_sums(4)(331) <= estimated(837) xor estimated(839);
partial_sums(4)(332) <= estimated(197) xor estimated(199);
partial_sums(4)(333) <= estimated(709) xor estimated(711);
partial_sums(4)(334) <= estimated(453) xor estimated(455);
partial_sums(4)(335) <= estimated(965) xor estimated(967);
partial_sums(4)(336) <= estimated(37) xor estimated(39);
partial_sums(4)(337) <= estimated(549) xor estimated(551);
partial_sums(4)(338) <= estimated(293) xor estimated(295);
partial_sums(4)(339) <= estimated(805) xor estimated(807);
partial_sums(4)(340) <= estimated(165) xor estimated(167);
partial_sums(4)(341) <= estimated(677) xor estimated(679);
partial_sums(4)(342) <= estimated(421) xor estimated(423);
partial_sums(4)(343) <= estimated(933) xor estimated(935);
partial_sums(4)(344) <= estimated(101) xor estimated(103);
partial_sums(4)(345) <= estimated(613) xor estimated(615);
partial_sums(4)(346) <= estimated(357) xor estimated(359);
partial_sums(4)(347) <= estimated(869) xor estimated(871);
partial_sums(4)(348) <= estimated(229) xor estimated(231);
partial_sums(4)(349) <= estimated(741) xor estimated(743);
partial_sums(4)(350) <= estimated(485) xor estimated(487);
partial_sums(4)(351) <= estimated(997) xor estimated(999);
partial_sums(4)(352) <= estimated(21) xor estimated(23);
partial_sums(4)(353) <= estimated(533) xor estimated(535);
partial_sums(4)(354) <= estimated(277) xor estimated(279);
partial_sums(4)(355) <= estimated(789) xor estimated(791);
partial_sums(4)(356) <= estimated(149) xor estimated(151);
partial_sums(4)(357) <= estimated(661) xor estimated(663);
partial_sums(4)(358) <= estimated(405) xor estimated(407);
partial_sums(4)(359) <= estimated(917) xor estimated(919);
partial_sums(4)(360) <= estimated(85) xor estimated(87);
partial_sums(4)(361) <= estimated(597) xor estimated(599);
partial_sums(4)(362) <= estimated(341) xor estimated(343);
partial_sums(4)(363) <= estimated(853) xor estimated(855);
partial_sums(4)(364) <= estimated(213) xor estimated(215);
partial_sums(4)(365) <= estimated(725) xor estimated(727);
partial_sums(4)(366) <= estimated(469) xor estimated(471);
partial_sums(4)(367) <= estimated(981) xor estimated(983);
partial_sums(4)(368) <= estimated(53) xor estimated(55);
partial_sums(4)(369) <= estimated(565) xor estimated(567);
partial_sums(4)(370) <= estimated(309) xor estimated(311);
partial_sums(4)(371) <= estimated(821) xor estimated(823);
partial_sums(4)(372) <= estimated(181) xor estimated(183);
partial_sums(4)(373) <= estimated(693) xor estimated(695);
partial_sums(4)(374) <= estimated(437) xor estimated(439);
partial_sums(4)(375) <= estimated(949) xor estimated(951);
partial_sums(4)(376) <= estimated(117) xor estimated(119);
partial_sums(4)(377) <= estimated(629) xor estimated(631);
partial_sums(4)(378) <= estimated(373) xor estimated(375);
partial_sums(4)(379) <= estimated(885) xor estimated(887);
partial_sums(4)(380) <= estimated(245) xor estimated(247);
partial_sums(4)(381) <= estimated(757) xor estimated(759);
partial_sums(4)(382) <= estimated(501) xor estimated(503);
partial_sums(4)(383) <= estimated(1013) xor estimated(1015);
partial_sums(4)(384) <= estimated(3) xor estimated(7);
partial_sums(4)(385) <= estimated(515) xor estimated(519);
partial_sums(4)(386) <= estimated(259) xor estimated(263);
partial_sums(4)(387) <= estimated(771) xor estimated(775);
partial_sums(4)(388) <= estimated(131) xor estimated(135);
partial_sums(4)(389) <= estimated(643) xor estimated(647);
partial_sums(4)(390) <= estimated(387) xor estimated(391);
partial_sums(4)(391) <= estimated(899) xor estimated(903);
partial_sums(4)(392) <= estimated(67) xor estimated(71);
partial_sums(4)(393) <= estimated(579) xor estimated(583);
partial_sums(4)(394) <= estimated(323) xor estimated(327);
partial_sums(4)(395) <= estimated(835) xor estimated(839);
partial_sums(4)(396) <= estimated(195) xor estimated(199);
partial_sums(4)(397) <= estimated(707) xor estimated(711);
partial_sums(4)(398) <= estimated(451) xor estimated(455);
partial_sums(4)(399) <= estimated(963) xor estimated(967);
partial_sums(4)(400) <= estimated(35) xor estimated(39);
partial_sums(4)(401) <= estimated(547) xor estimated(551);
partial_sums(4)(402) <= estimated(291) xor estimated(295);
partial_sums(4)(403) <= estimated(803) xor estimated(807);
partial_sums(4)(404) <= estimated(163) xor estimated(167);
partial_sums(4)(405) <= estimated(675) xor estimated(679);
partial_sums(4)(406) <= estimated(419) xor estimated(423);
partial_sums(4)(407) <= estimated(931) xor estimated(935);
partial_sums(4)(408) <= estimated(99) xor estimated(103);
partial_sums(4)(409) <= estimated(611) xor estimated(615);
partial_sums(4)(410) <= estimated(355) xor estimated(359);
partial_sums(4)(411) <= estimated(867) xor estimated(871);
partial_sums(4)(412) <= estimated(227) xor estimated(231);
partial_sums(4)(413) <= estimated(739) xor estimated(743);
partial_sums(4)(414) <= estimated(483) xor estimated(487);
partial_sums(4)(415) <= estimated(995) xor estimated(999);
partial_sums(4)(416) <= estimated(19) xor estimated(23);
partial_sums(4)(417) <= estimated(531) xor estimated(535);
partial_sums(4)(418) <= estimated(275) xor estimated(279);
partial_sums(4)(419) <= estimated(787) xor estimated(791);
partial_sums(4)(420) <= estimated(147) xor estimated(151);
partial_sums(4)(421) <= estimated(659) xor estimated(663);
partial_sums(4)(422) <= estimated(403) xor estimated(407);
partial_sums(4)(423) <= estimated(915) xor estimated(919);
partial_sums(4)(424) <= estimated(83) xor estimated(87);
partial_sums(4)(425) <= estimated(595) xor estimated(599);
partial_sums(4)(426) <= estimated(339) xor estimated(343);
partial_sums(4)(427) <= estimated(851) xor estimated(855);
partial_sums(4)(428) <= estimated(211) xor estimated(215);
partial_sums(4)(429) <= estimated(723) xor estimated(727);
partial_sums(4)(430) <= estimated(467) xor estimated(471);
partial_sums(4)(431) <= estimated(979) xor estimated(983);
partial_sums(4)(432) <= estimated(51) xor estimated(55);
partial_sums(4)(433) <= estimated(563) xor estimated(567);
partial_sums(4)(434) <= estimated(307) xor estimated(311);
partial_sums(4)(435) <= estimated(819) xor estimated(823);
partial_sums(4)(436) <= estimated(179) xor estimated(183);
partial_sums(4)(437) <= estimated(691) xor estimated(695);
partial_sums(4)(438) <= estimated(435) xor estimated(439);
partial_sums(4)(439) <= estimated(947) xor estimated(951);
partial_sums(4)(440) <= estimated(115) xor estimated(119);
partial_sums(4)(441) <= estimated(627) xor estimated(631);
partial_sums(4)(442) <= estimated(371) xor estimated(375);
partial_sums(4)(443) <= estimated(883) xor estimated(887);
partial_sums(4)(444) <= estimated(243) xor estimated(247);
partial_sums(4)(445) <= estimated(755) xor estimated(759);
partial_sums(4)(446) <= estimated(499) xor estimated(503);
partial_sums(4)(447) <= estimated(1011) xor estimated(1015);
partial_sums(4)(448) <= estimated(7);
partial_sums(4)(449) <= estimated(519);
partial_sums(4)(450) <= estimated(263);
partial_sums(4)(451) <= estimated(775);
partial_sums(4)(452) <= estimated(135);
partial_sums(4)(453) <= estimated(647);
partial_sums(4)(454) <= estimated(391);
partial_sums(4)(455) <= estimated(903);
partial_sums(4)(456) <= estimated(71);
partial_sums(4)(457) <= estimated(583);
partial_sums(4)(458) <= estimated(327);
partial_sums(4)(459) <= estimated(839);
partial_sums(4)(460) <= estimated(199);
partial_sums(4)(461) <= estimated(711);
partial_sums(4)(462) <= estimated(455);
partial_sums(4)(463) <= estimated(967);
partial_sums(4)(464) <= estimated(39);
partial_sums(4)(465) <= estimated(551);
partial_sums(4)(466) <= estimated(295);
partial_sums(4)(467) <= estimated(807);
partial_sums(4)(468) <= estimated(167);
partial_sums(4)(469) <= estimated(679);
partial_sums(4)(470) <= estimated(423);
partial_sums(4)(471) <= estimated(935);
partial_sums(4)(472) <= estimated(103);
partial_sums(4)(473) <= estimated(615);
partial_sums(4)(474) <= estimated(359);
partial_sums(4)(475) <= estimated(871);
partial_sums(4)(476) <= estimated(231);
partial_sums(4)(477) <= estimated(743);
partial_sums(4)(478) <= estimated(487);
partial_sums(4)(479) <= estimated(999);
partial_sums(4)(480) <= estimated(23);
partial_sums(4)(481) <= estimated(535);
partial_sums(4)(482) <= estimated(279);
partial_sums(4)(483) <= estimated(791);
partial_sums(4)(484) <= estimated(151);
partial_sums(4)(485) <= estimated(663);
partial_sums(4)(486) <= estimated(407);
partial_sums(4)(487) <= estimated(919);
partial_sums(4)(488) <= estimated(87);
partial_sums(4)(489) <= estimated(599);
partial_sums(4)(490) <= estimated(343);
partial_sums(4)(491) <= estimated(855);
partial_sums(4)(492) <= estimated(215);
partial_sums(4)(493) <= estimated(727);
partial_sums(4)(494) <= estimated(471);
partial_sums(4)(495) <= estimated(983);
partial_sums(4)(496) <= estimated(55);
partial_sums(4)(497) <= estimated(567);
partial_sums(4)(498) <= estimated(311);
partial_sums(4)(499) <= estimated(823);
partial_sums(4)(500) <= estimated(183);
partial_sums(4)(501) <= estimated(695);
partial_sums(4)(502) <= estimated(439);
partial_sums(4)(503) <= estimated(951);
partial_sums(4)(504) <= estimated(119);
partial_sums(4)(505) <= estimated(631);
partial_sums(4)(506) <= estimated(375);
partial_sums(4)(507) <= estimated(887);
partial_sums(4)(508) <= estimated(247);
partial_sums(4)(509) <= estimated(759);
partial_sums(4)(510) <= estimated(503);
partial_sums(4)(511) <= estimated(1015);
partial_sums(5)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(1) <= estimated(512) xor estimated(513) xor estimated(514) xor estimated(515) xor estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527);
partial_sums(5)(2) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(3) <= estimated(768) xor estimated(769) xor estimated(770) xor estimated(771) xor estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783);
partial_sums(5)(4) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(5) <= estimated(640) xor estimated(641) xor estimated(642) xor estimated(643) xor estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655);
partial_sums(5)(6) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(7) <= estimated(896) xor estimated(897) xor estimated(898) xor estimated(899) xor estimated(900) xor estimated(901) xor estimated(902) xor estimated(903) xor estimated(904) xor estimated(905) xor estimated(906) xor estimated(907) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911);
partial_sums(5)(8) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(9) <= estimated(576) xor estimated(577) xor estimated(578) xor estimated(579) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591);
partial_sums(5)(10) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(11) <= estimated(832) xor estimated(833) xor estimated(834) xor estimated(835) xor estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847);
partial_sums(5)(12) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(13) <= estimated(704) xor estimated(705) xor estimated(706) xor estimated(707) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719);
partial_sums(5)(14) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(15) <= estimated(960) xor estimated(961) xor estimated(962) xor estimated(963) xor estimated(964) xor estimated(965) xor estimated(966) xor estimated(967) xor estimated(968) xor estimated(969) xor estimated(970) xor estimated(971) xor estimated(972) xor estimated(973) xor estimated(974) xor estimated(975);
partial_sums(5)(16) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(17) <= estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559);
partial_sums(5)(18) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(19) <= estimated(800) xor estimated(801) xor estimated(802) xor estimated(803) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815);
partial_sums(5)(20) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(21) <= estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687);
partial_sums(5)(22) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(23) <= estimated(928) xor estimated(929) xor estimated(930) xor estimated(931) xor estimated(932) xor estimated(933) xor estimated(934) xor estimated(935) xor estimated(936) xor estimated(937) xor estimated(938) xor estimated(939) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943);
partial_sums(5)(24) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(25) <= estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623);
partial_sums(5)(26) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(27) <= estimated(864) xor estimated(865) xor estimated(866) xor estimated(867) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879);
partial_sums(5)(28) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(29) <= estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751);
partial_sums(5)(30) <= estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(31) <= estimated(992) xor estimated(993) xor estimated(994) xor estimated(995) xor estimated(996) xor estimated(997) xor estimated(998) xor estimated(999) xor estimated(1000) xor estimated(1001) xor estimated(1002) xor estimated(1003) xor estimated(1004) xor estimated(1005) xor estimated(1006) xor estimated(1007);
partial_sums(5)(32) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(33) <= estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527);
partial_sums(5)(34) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(35) <= estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783);
partial_sums(5)(36) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(37) <= estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655);
partial_sums(5)(38) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(39) <= estimated(904) xor estimated(905) xor estimated(906) xor estimated(907) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911);
partial_sums(5)(40) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(41) <= estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591);
partial_sums(5)(42) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(43) <= estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847);
partial_sums(5)(44) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(45) <= estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719);
partial_sums(5)(46) <= estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(47) <= estimated(968) xor estimated(969) xor estimated(970) xor estimated(971) xor estimated(972) xor estimated(973) xor estimated(974) xor estimated(975);
partial_sums(5)(48) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(49) <= estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559);
partial_sums(5)(50) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(51) <= estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815);
partial_sums(5)(52) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(53) <= estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687);
partial_sums(5)(54) <= estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(55) <= estimated(936) xor estimated(937) xor estimated(938) xor estimated(939) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943);
partial_sums(5)(56) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(57) <= estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623);
partial_sums(5)(58) <= estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(59) <= estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879);
partial_sums(5)(60) <= estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(61) <= estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751);
partial_sums(5)(62) <= estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(63) <= estimated(1000) xor estimated(1001) xor estimated(1002) xor estimated(1003) xor estimated(1004) xor estimated(1005) xor estimated(1006) xor estimated(1007);
partial_sums(5)(64) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(65) <= estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527);
partial_sums(5)(66) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(67) <= estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783);
partial_sums(5)(68) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(69) <= estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655);
partial_sums(5)(70) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(71) <= estimated(900) xor estimated(901) xor estimated(902) xor estimated(903) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911);
partial_sums(5)(72) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(73) <= estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591);
partial_sums(5)(74) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(75) <= estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847);
partial_sums(5)(76) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(77) <= estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719);
partial_sums(5)(78) <= estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(79) <= estimated(964) xor estimated(965) xor estimated(966) xor estimated(967) xor estimated(972) xor estimated(973) xor estimated(974) xor estimated(975);
partial_sums(5)(80) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(81) <= estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559);
partial_sums(5)(82) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(83) <= estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815);
partial_sums(5)(84) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(85) <= estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687);
partial_sums(5)(86) <= estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(87) <= estimated(932) xor estimated(933) xor estimated(934) xor estimated(935) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943);
partial_sums(5)(88) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(89) <= estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623);
partial_sums(5)(90) <= estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(91) <= estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879);
partial_sums(5)(92) <= estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(93) <= estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751);
partial_sums(5)(94) <= estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(95) <= estimated(996) xor estimated(997) xor estimated(998) xor estimated(999) xor estimated(1004) xor estimated(1005) xor estimated(1006) xor estimated(1007);
partial_sums(5)(96) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15);
partial_sums(5)(97) <= estimated(524) xor estimated(525) xor estimated(526) xor estimated(527);
partial_sums(5)(98) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271);
partial_sums(5)(99) <= estimated(780) xor estimated(781) xor estimated(782) xor estimated(783);
partial_sums(5)(100) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143);
partial_sums(5)(101) <= estimated(652) xor estimated(653) xor estimated(654) xor estimated(655);
partial_sums(5)(102) <= estimated(396) xor estimated(397) xor estimated(398) xor estimated(399);
partial_sums(5)(103) <= estimated(908) xor estimated(909) xor estimated(910) xor estimated(911);
partial_sums(5)(104) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79);
partial_sums(5)(105) <= estimated(588) xor estimated(589) xor estimated(590) xor estimated(591);
partial_sums(5)(106) <= estimated(332) xor estimated(333) xor estimated(334) xor estimated(335);
partial_sums(5)(107) <= estimated(844) xor estimated(845) xor estimated(846) xor estimated(847);
partial_sums(5)(108) <= estimated(204) xor estimated(205) xor estimated(206) xor estimated(207);
partial_sums(5)(109) <= estimated(716) xor estimated(717) xor estimated(718) xor estimated(719);
partial_sums(5)(110) <= estimated(460) xor estimated(461) xor estimated(462) xor estimated(463);
partial_sums(5)(111) <= estimated(972) xor estimated(973) xor estimated(974) xor estimated(975);
partial_sums(5)(112) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47);
partial_sums(5)(113) <= estimated(556) xor estimated(557) xor estimated(558) xor estimated(559);
partial_sums(5)(114) <= estimated(300) xor estimated(301) xor estimated(302) xor estimated(303);
partial_sums(5)(115) <= estimated(812) xor estimated(813) xor estimated(814) xor estimated(815);
partial_sums(5)(116) <= estimated(172) xor estimated(173) xor estimated(174) xor estimated(175);
partial_sums(5)(117) <= estimated(684) xor estimated(685) xor estimated(686) xor estimated(687);
partial_sums(5)(118) <= estimated(428) xor estimated(429) xor estimated(430) xor estimated(431);
partial_sums(5)(119) <= estimated(940) xor estimated(941) xor estimated(942) xor estimated(943);
partial_sums(5)(120) <= estimated(108) xor estimated(109) xor estimated(110) xor estimated(111);
partial_sums(5)(121) <= estimated(620) xor estimated(621) xor estimated(622) xor estimated(623);
partial_sums(5)(122) <= estimated(364) xor estimated(365) xor estimated(366) xor estimated(367);
partial_sums(5)(123) <= estimated(876) xor estimated(877) xor estimated(878) xor estimated(879);
partial_sums(5)(124) <= estimated(236) xor estimated(237) xor estimated(238) xor estimated(239);
partial_sums(5)(125) <= estimated(748) xor estimated(749) xor estimated(750) xor estimated(751);
partial_sums(5)(126) <= estimated(492) xor estimated(493) xor estimated(494) xor estimated(495);
partial_sums(5)(127) <= estimated(1004) xor estimated(1005) xor estimated(1006) xor estimated(1007);
partial_sums(5)(128) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15);
partial_sums(5)(129) <= estimated(514) xor estimated(515) xor estimated(518) xor estimated(519) xor estimated(522) xor estimated(523) xor estimated(526) xor estimated(527);
partial_sums(5)(130) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271);
partial_sums(5)(131) <= estimated(770) xor estimated(771) xor estimated(774) xor estimated(775) xor estimated(778) xor estimated(779) xor estimated(782) xor estimated(783);
partial_sums(5)(132) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143);
partial_sums(5)(133) <= estimated(642) xor estimated(643) xor estimated(646) xor estimated(647) xor estimated(650) xor estimated(651) xor estimated(654) xor estimated(655);
partial_sums(5)(134) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399);
partial_sums(5)(135) <= estimated(898) xor estimated(899) xor estimated(902) xor estimated(903) xor estimated(906) xor estimated(907) xor estimated(910) xor estimated(911);
partial_sums(5)(136) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79);
partial_sums(5)(137) <= estimated(578) xor estimated(579) xor estimated(582) xor estimated(583) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591);
partial_sums(5)(138) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335);
partial_sums(5)(139) <= estimated(834) xor estimated(835) xor estimated(838) xor estimated(839) xor estimated(842) xor estimated(843) xor estimated(846) xor estimated(847);
partial_sums(5)(140) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207);
partial_sums(5)(141) <= estimated(706) xor estimated(707) xor estimated(710) xor estimated(711) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719);
partial_sums(5)(142) <= estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463);
partial_sums(5)(143) <= estimated(962) xor estimated(963) xor estimated(966) xor estimated(967) xor estimated(970) xor estimated(971) xor estimated(974) xor estimated(975);
partial_sums(5)(144) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47);
partial_sums(5)(145) <= estimated(546) xor estimated(547) xor estimated(550) xor estimated(551) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559);
partial_sums(5)(146) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303);
partial_sums(5)(147) <= estimated(802) xor estimated(803) xor estimated(806) xor estimated(807) xor estimated(810) xor estimated(811) xor estimated(814) xor estimated(815);
partial_sums(5)(148) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175);
partial_sums(5)(149) <= estimated(674) xor estimated(675) xor estimated(678) xor estimated(679) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687);
partial_sums(5)(150) <= estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431);
partial_sums(5)(151) <= estimated(930) xor estimated(931) xor estimated(934) xor estimated(935) xor estimated(938) xor estimated(939) xor estimated(942) xor estimated(943);
partial_sums(5)(152) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111);
partial_sums(5)(153) <= estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623);
partial_sums(5)(154) <= estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367);
partial_sums(5)(155) <= estimated(866) xor estimated(867) xor estimated(870) xor estimated(871) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879);
partial_sums(5)(156) <= estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239);
partial_sums(5)(157) <= estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751);
partial_sums(5)(158) <= estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495);
partial_sums(5)(159) <= estimated(994) xor estimated(995) xor estimated(998) xor estimated(999) xor estimated(1002) xor estimated(1003) xor estimated(1006) xor estimated(1007);
partial_sums(5)(160) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15);
partial_sums(5)(161) <= estimated(522) xor estimated(523) xor estimated(526) xor estimated(527);
partial_sums(5)(162) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271);
partial_sums(5)(163) <= estimated(778) xor estimated(779) xor estimated(782) xor estimated(783);
partial_sums(5)(164) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143);
partial_sums(5)(165) <= estimated(650) xor estimated(651) xor estimated(654) xor estimated(655);
partial_sums(5)(166) <= estimated(394) xor estimated(395) xor estimated(398) xor estimated(399);
partial_sums(5)(167) <= estimated(906) xor estimated(907) xor estimated(910) xor estimated(911);
partial_sums(5)(168) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79);
partial_sums(5)(169) <= estimated(586) xor estimated(587) xor estimated(590) xor estimated(591);
partial_sums(5)(170) <= estimated(330) xor estimated(331) xor estimated(334) xor estimated(335);
partial_sums(5)(171) <= estimated(842) xor estimated(843) xor estimated(846) xor estimated(847);
partial_sums(5)(172) <= estimated(202) xor estimated(203) xor estimated(206) xor estimated(207);
partial_sums(5)(173) <= estimated(714) xor estimated(715) xor estimated(718) xor estimated(719);
partial_sums(5)(174) <= estimated(458) xor estimated(459) xor estimated(462) xor estimated(463);
partial_sums(5)(175) <= estimated(970) xor estimated(971) xor estimated(974) xor estimated(975);
partial_sums(5)(176) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47);
partial_sums(5)(177) <= estimated(554) xor estimated(555) xor estimated(558) xor estimated(559);
partial_sums(5)(178) <= estimated(298) xor estimated(299) xor estimated(302) xor estimated(303);
partial_sums(5)(179) <= estimated(810) xor estimated(811) xor estimated(814) xor estimated(815);
partial_sums(5)(180) <= estimated(170) xor estimated(171) xor estimated(174) xor estimated(175);
partial_sums(5)(181) <= estimated(682) xor estimated(683) xor estimated(686) xor estimated(687);
partial_sums(5)(182) <= estimated(426) xor estimated(427) xor estimated(430) xor estimated(431);
partial_sums(5)(183) <= estimated(938) xor estimated(939) xor estimated(942) xor estimated(943);
partial_sums(5)(184) <= estimated(106) xor estimated(107) xor estimated(110) xor estimated(111);
partial_sums(5)(185) <= estimated(618) xor estimated(619) xor estimated(622) xor estimated(623);
partial_sums(5)(186) <= estimated(362) xor estimated(363) xor estimated(366) xor estimated(367);
partial_sums(5)(187) <= estimated(874) xor estimated(875) xor estimated(878) xor estimated(879);
partial_sums(5)(188) <= estimated(234) xor estimated(235) xor estimated(238) xor estimated(239);
partial_sums(5)(189) <= estimated(746) xor estimated(747) xor estimated(750) xor estimated(751);
partial_sums(5)(190) <= estimated(490) xor estimated(491) xor estimated(494) xor estimated(495);
partial_sums(5)(191) <= estimated(1002) xor estimated(1003) xor estimated(1006) xor estimated(1007);
partial_sums(5)(192) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15);
partial_sums(5)(193) <= estimated(518) xor estimated(519) xor estimated(526) xor estimated(527);
partial_sums(5)(194) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271);
partial_sums(5)(195) <= estimated(774) xor estimated(775) xor estimated(782) xor estimated(783);
partial_sums(5)(196) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143);
partial_sums(5)(197) <= estimated(646) xor estimated(647) xor estimated(654) xor estimated(655);
partial_sums(5)(198) <= estimated(390) xor estimated(391) xor estimated(398) xor estimated(399);
partial_sums(5)(199) <= estimated(902) xor estimated(903) xor estimated(910) xor estimated(911);
partial_sums(5)(200) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79);
partial_sums(5)(201) <= estimated(582) xor estimated(583) xor estimated(590) xor estimated(591);
partial_sums(5)(202) <= estimated(326) xor estimated(327) xor estimated(334) xor estimated(335);
partial_sums(5)(203) <= estimated(838) xor estimated(839) xor estimated(846) xor estimated(847);
partial_sums(5)(204) <= estimated(198) xor estimated(199) xor estimated(206) xor estimated(207);
partial_sums(5)(205) <= estimated(710) xor estimated(711) xor estimated(718) xor estimated(719);
partial_sums(5)(206) <= estimated(454) xor estimated(455) xor estimated(462) xor estimated(463);
partial_sums(5)(207) <= estimated(966) xor estimated(967) xor estimated(974) xor estimated(975);
partial_sums(5)(208) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47);
partial_sums(5)(209) <= estimated(550) xor estimated(551) xor estimated(558) xor estimated(559);
partial_sums(5)(210) <= estimated(294) xor estimated(295) xor estimated(302) xor estimated(303);
partial_sums(5)(211) <= estimated(806) xor estimated(807) xor estimated(814) xor estimated(815);
partial_sums(5)(212) <= estimated(166) xor estimated(167) xor estimated(174) xor estimated(175);
partial_sums(5)(213) <= estimated(678) xor estimated(679) xor estimated(686) xor estimated(687);
partial_sums(5)(214) <= estimated(422) xor estimated(423) xor estimated(430) xor estimated(431);
partial_sums(5)(215) <= estimated(934) xor estimated(935) xor estimated(942) xor estimated(943);
partial_sums(5)(216) <= estimated(102) xor estimated(103) xor estimated(110) xor estimated(111);
partial_sums(5)(217) <= estimated(614) xor estimated(615) xor estimated(622) xor estimated(623);
partial_sums(5)(218) <= estimated(358) xor estimated(359) xor estimated(366) xor estimated(367);
partial_sums(5)(219) <= estimated(870) xor estimated(871) xor estimated(878) xor estimated(879);
partial_sums(5)(220) <= estimated(230) xor estimated(231) xor estimated(238) xor estimated(239);
partial_sums(5)(221) <= estimated(742) xor estimated(743) xor estimated(750) xor estimated(751);
partial_sums(5)(222) <= estimated(486) xor estimated(487) xor estimated(494) xor estimated(495);
partial_sums(5)(223) <= estimated(998) xor estimated(999) xor estimated(1006) xor estimated(1007);
partial_sums(5)(224) <= estimated(14) xor estimated(15);
partial_sums(5)(225) <= estimated(526) xor estimated(527);
partial_sums(5)(226) <= estimated(270) xor estimated(271);
partial_sums(5)(227) <= estimated(782) xor estimated(783);
partial_sums(5)(228) <= estimated(142) xor estimated(143);
partial_sums(5)(229) <= estimated(654) xor estimated(655);
partial_sums(5)(230) <= estimated(398) xor estimated(399);
partial_sums(5)(231) <= estimated(910) xor estimated(911);
partial_sums(5)(232) <= estimated(78) xor estimated(79);
partial_sums(5)(233) <= estimated(590) xor estimated(591);
partial_sums(5)(234) <= estimated(334) xor estimated(335);
partial_sums(5)(235) <= estimated(846) xor estimated(847);
partial_sums(5)(236) <= estimated(206) xor estimated(207);
partial_sums(5)(237) <= estimated(718) xor estimated(719);
partial_sums(5)(238) <= estimated(462) xor estimated(463);
partial_sums(5)(239) <= estimated(974) xor estimated(975);
partial_sums(5)(240) <= estimated(46) xor estimated(47);
partial_sums(5)(241) <= estimated(558) xor estimated(559);
partial_sums(5)(242) <= estimated(302) xor estimated(303);
partial_sums(5)(243) <= estimated(814) xor estimated(815);
partial_sums(5)(244) <= estimated(174) xor estimated(175);
partial_sums(5)(245) <= estimated(686) xor estimated(687);
partial_sums(5)(246) <= estimated(430) xor estimated(431);
partial_sums(5)(247) <= estimated(942) xor estimated(943);
partial_sums(5)(248) <= estimated(110) xor estimated(111);
partial_sums(5)(249) <= estimated(622) xor estimated(623);
partial_sums(5)(250) <= estimated(366) xor estimated(367);
partial_sums(5)(251) <= estimated(878) xor estimated(879);
partial_sums(5)(252) <= estimated(238) xor estimated(239);
partial_sums(5)(253) <= estimated(750) xor estimated(751);
partial_sums(5)(254) <= estimated(494) xor estimated(495);
partial_sums(5)(255) <= estimated(1006) xor estimated(1007);
partial_sums(5)(256) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15);
partial_sums(5)(257) <= estimated(513) xor estimated(515) xor estimated(517) xor estimated(519) xor estimated(521) xor estimated(523) xor estimated(525) xor estimated(527);
partial_sums(5)(258) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271);
partial_sums(5)(259) <= estimated(769) xor estimated(771) xor estimated(773) xor estimated(775) xor estimated(777) xor estimated(779) xor estimated(781) xor estimated(783);
partial_sums(5)(260) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143);
partial_sums(5)(261) <= estimated(641) xor estimated(643) xor estimated(645) xor estimated(647) xor estimated(649) xor estimated(651) xor estimated(653) xor estimated(655);
partial_sums(5)(262) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399);
partial_sums(5)(263) <= estimated(897) xor estimated(899) xor estimated(901) xor estimated(903) xor estimated(905) xor estimated(907) xor estimated(909) xor estimated(911);
partial_sums(5)(264) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79);
partial_sums(5)(265) <= estimated(577) xor estimated(579) xor estimated(581) xor estimated(583) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591);
partial_sums(5)(266) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335);
partial_sums(5)(267) <= estimated(833) xor estimated(835) xor estimated(837) xor estimated(839) xor estimated(841) xor estimated(843) xor estimated(845) xor estimated(847);
partial_sums(5)(268) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207);
partial_sums(5)(269) <= estimated(705) xor estimated(707) xor estimated(709) xor estimated(711) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719);
partial_sums(5)(270) <= estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463);
partial_sums(5)(271) <= estimated(961) xor estimated(963) xor estimated(965) xor estimated(967) xor estimated(969) xor estimated(971) xor estimated(973) xor estimated(975);
partial_sums(5)(272) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47);
partial_sums(5)(273) <= estimated(545) xor estimated(547) xor estimated(549) xor estimated(551) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559);
partial_sums(5)(274) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303);
partial_sums(5)(275) <= estimated(801) xor estimated(803) xor estimated(805) xor estimated(807) xor estimated(809) xor estimated(811) xor estimated(813) xor estimated(815);
partial_sums(5)(276) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175);
partial_sums(5)(277) <= estimated(673) xor estimated(675) xor estimated(677) xor estimated(679) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687);
partial_sums(5)(278) <= estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431);
partial_sums(5)(279) <= estimated(929) xor estimated(931) xor estimated(933) xor estimated(935) xor estimated(937) xor estimated(939) xor estimated(941) xor estimated(943);
partial_sums(5)(280) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111);
partial_sums(5)(281) <= estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623);
partial_sums(5)(282) <= estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367);
partial_sums(5)(283) <= estimated(865) xor estimated(867) xor estimated(869) xor estimated(871) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879);
partial_sums(5)(284) <= estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239);
partial_sums(5)(285) <= estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751);
partial_sums(5)(286) <= estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495);
partial_sums(5)(287) <= estimated(993) xor estimated(995) xor estimated(997) xor estimated(999) xor estimated(1001) xor estimated(1003) xor estimated(1005) xor estimated(1007);
partial_sums(5)(288) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15);
partial_sums(5)(289) <= estimated(521) xor estimated(523) xor estimated(525) xor estimated(527);
partial_sums(5)(290) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271);
partial_sums(5)(291) <= estimated(777) xor estimated(779) xor estimated(781) xor estimated(783);
partial_sums(5)(292) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143);
partial_sums(5)(293) <= estimated(649) xor estimated(651) xor estimated(653) xor estimated(655);
partial_sums(5)(294) <= estimated(393) xor estimated(395) xor estimated(397) xor estimated(399);
partial_sums(5)(295) <= estimated(905) xor estimated(907) xor estimated(909) xor estimated(911);
partial_sums(5)(296) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79);
partial_sums(5)(297) <= estimated(585) xor estimated(587) xor estimated(589) xor estimated(591);
partial_sums(5)(298) <= estimated(329) xor estimated(331) xor estimated(333) xor estimated(335);
partial_sums(5)(299) <= estimated(841) xor estimated(843) xor estimated(845) xor estimated(847);
partial_sums(5)(300) <= estimated(201) xor estimated(203) xor estimated(205) xor estimated(207);
partial_sums(5)(301) <= estimated(713) xor estimated(715) xor estimated(717) xor estimated(719);
partial_sums(5)(302) <= estimated(457) xor estimated(459) xor estimated(461) xor estimated(463);
partial_sums(5)(303) <= estimated(969) xor estimated(971) xor estimated(973) xor estimated(975);
partial_sums(5)(304) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47);
partial_sums(5)(305) <= estimated(553) xor estimated(555) xor estimated(557) xor estimated(559);
partial_sums(5)(306) <= estimated(297) xor estimated(299) xor estimated(301) xor estimated(303);
partial_sums(5)(307) <= estimated(809) xor estimated(811) xor estimated(813) xor estimated(815);
partial_sums(5)(308) <= estimated(169) xor estimated(171) xor estimated(173) xor estimated(175);
partial_sums(5)(309) <= estimated(681) xor estimated(683) xor estimated(685) xor estimated(687);
partial_sums(5)(310) <= estimated(425) xor estimated(427) xor estimated(429) xor estimated(431);
partial_sums(5)(311) <= estimated(937) xor estimated(939) xor estimated(941) xor estimated(943);
partial_sums(5)(312) <= estimated(105) xor estimated(107) xor estimated(109) xor estimated(111);
partial_sums(5)(313) <= estimated(617) xor estimated(619) xor estimated(621) xor estimated(623);
partial_sums(5)(314) <= estimated(361) xor estimated(363) xor estimated(365) xor estimated(367);
partial_sums(5)(315) <= estimated(873) xor estimated(875) xor estimated(877) xor estimated(879);
partial_sums(5)(316) <= estimated(233) xor estimated(235) xor estimated(237) xor estimated(239);
partial_sums(5)(317) <= estimated(745) xor estimated(747) xor estimated(749) xor estimated(751);
partial_sums(5)(318) <= estimated(489) xor estimated(491) xor estimated(493) xor estimated(495);
partial_sums(5)(319) <= estimated(1001) xor estimated(1003) xor estimated(1005) xor estimated(1007);
partial_sums(5)(320) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15);
partial_sums(5)(321) <= estimated(517) xor estimated(519) xor estimated(525) xor estimated(527);
partial_sums(5)(322) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271);
partial_sums(5)(323) <= estimated(773) xor estimated(775) xor estimated(781) xor estimated(783);
partial_sums(5)(324) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143);
partial_sums(5)(325) <= estimated(645) xor estimated(647) xor estimated(653) xor estimated(655);
partial_sums(5)(326) <= estimated(389) xor estimated(391) xor estimated(397) xor estimated(399);
partial_sums(5)(327) <= estimated(901) xor estimated(903) xor estimated(909) xor estimated(911);
partial_sums(5)(328) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79);
partial_sums(5)(329) <= estimated(581) xor estimated(583) xor estimated(589) xor estimated(591);
partial_sums(5)(330) <= estimated(325) xor estimated(327) xor estimated(333) xor estimated(335);
partial_sums(5)(331) <= estimated(837) xor estimated(839) xor estimated(845) xor estimated(847);
partial_sums(5)(332) <= estimated(197) xor estimated(199) xor estimated(205) xor estimated(207);
partial_sums(5)(333) <= estimated(709) xor estimated(711) xor estimated(717) xor estimated(719);
partial_sums(5)(334) <= estimated(453) xor estimated(455) xor estimated(461) xor estimated(463);
partial_sums(5)(335) <= estimated(965) xor estimated(967) xor estimated(973) xor estimated(975);
partial_sums(5)(336) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47);
partial_sums(5)(337) <= estimated(549) xor estimated(551) xor estimated(557) xor estimated(559);
partial_sums(5)(338) <= estimated(293) xor estimated(295) xor estimated(301) xor estimated(303);
partial_sums(5)(339) <= estimated(805) xor estimated(807) xor estimated(813) xor estimated(815);
partial_sums(5)(340) <= estimated(165) xor estimated(167) xor estimated(173) xor estimated(175);
partial_sums(5)(341) <= estimated(677) xor estimated(679) xor estimated(685) xor estimated(687);
partial_sums(5)(342) <= estimated(421) xor estimated(423) xor estimated(429) xor estimated(431);
partial_sums(5)(343) <= estimated(933) xor estimated(935) xor estimated(941) xor estimated(943);
partial_sums(5)(344) <= estimated(101) xor estimated(103) xor estimated(109) xor estimated(111);
partial_sums(5)(345) <= estimated(613) xor estimated(615) xor estimated(621) xor estimated(623);
partial_sums(5)(346) <= estimated(357) xor estimated(359) xor estimated(365) xor estimated(367);
partial_sums(5)(347) <= estimated(869) xor estimated(871) xor estimated(877) xor estimated(879);
partial_sums(5)(348) <= estimated(229) xor estimated(231) xor estimated(237) xor estimated(239);
partial_sums(5)(349) <= estimated(741) xor estimated(743) xor estimated(749) xor estimated(751);
partial_sums(5)(350) <= estimated(485) xor estimated(487) xor estimated(493) xor estimated(495);
partial_sums(5)(351) <= estimated(997) xor estimated(999) xor estimated(1005) xor estimated(1007);
partial_sums(5)(352) <= estimated(13) xor estimated(15);
partial_sums(5)(353) <= estimated(525) xor estimated(527);
partial_sums(5)(354) <= estimated(269) xor estimated(271);
partial_sums(5)(355) <= estimated(781) xor estimated(783);
partial_sums(5)(356) <= estimated(141) xor estimated(143);
partial_sums(5)(357) <= estimated(653) xor estimated(655);
partial_sums(5)(358) <= estimated(397) xor estimated(399);
partial_sums(5)(359) <= estimated(909) xor estimated(911);
partial_sums(5)(360) <= estimated(77) xor estimated(79);
partial_sums(5)(361) <= estimated(589) xor estimated(591);
partial_sums(5)(362) <= estimated(333) xor estimated(335);
partial_sums(5)(363) <= estimated(845) xor estimated(847);
partial_sums(5)(364) <= estimated(205) xor estimated(207);
partial_sums(5)(365) <= estimated(717) xor estimated(719);
partial_sums(5)(366) <= estimated(461) xor estimated(463);
partial_sums(5)(367) <= estimated(973) xor estimated(975);
partial_sums(5)(368) <= estimated(45) xor estimated(47);
partial_sums(5)(369) <= estimated(557) xor estimated(559);
partial_sums(5)(370) <= estimated(301) xor estimated(303);
partial_sums(5)(371) <= estimated(813) xor estimated(815);
partial_sums(5)(372) <= estimated(173) xor estimated(175);
partial_sums(5)(373) <= estimated(685) xor estimated(687);
partial_sums(5)(374) <= estimated(429) xor estimated(431);
partial_sums(5)(375) <= estimated(941) xor estimated(943);
partial_sums(5)(376) <= estimated(109) xor estimated(111);
partial_sums(5)(377) <= estimated(621) xor estimated(623);
partial_sums(5)(378) <= estimated(365) xor estimated(367);
partial_sums(5)(379) <= estimated(877) xor estimated(879);
partial_sums(5)(380) <= estimated(237) xor estimated(239);
partial_sums(5)(381) <= estimated(749) xor estimated(751);
partial_sums(5)(382) <= estimated(493) xor estimated(495);
partial_sums(5)(383) <= estimated(1005) xor estimated(1007);
partial_sums(5)(384) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15);
partial_sums(5)(385) <= estimated(515) xor estimated(519) xor estimated(523) xor estimated(527);
partial_sums(5)(386) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271);
partial_sums(5)(387) <= estimated(771) xor estimated(775) xor estimated(779) xor estimated(783);
partial_sums(5)(388) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143);
partial_sums(5)(389) <= estimated(643) xor estimated(647) xor estimated(651) xor estimated(655);
partial_sums(5)(390) <= estimated(387) xor estimated(391) xor estimated(395) xor estimated(399);
partial_sums(5)(391) <= estimated(899) xor estimated(903) xor estimated(907) xor estimated(911);
partial_sums(5)(392) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79);
partial_sums(5)(393) <= estimated(579) xor estimated(583) xor estimated(587) xor estimated(591);
partial_sums(5)(394) <= estimated(323) xor estimated(327) xor estimated(331) xor estimated(335);
partial_sums(5)(395) <= estimated(835) xor estimated(839) xor estimated(843) xor estimated(847);
partial_sums(5)(396) <= estimated(195) xor estimated(199) xor estimated(203) xor estimated(207);
partial_sums(5)(397) <= estimated(707) xor estimated(711) xor estimated(715) xor estimated(719);
partial_sums(5)(398) <= estimated(451) xor estimated(455) xor estimated(459) xor estimated(463);
partial_sums(5)(399) <= estimated(963) xor estimated(967) xor estimated(971) xor estimated(975);
partial_sums(5)(400) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47);
partial_sums(5)(401) <= estimated(547) xor estimated(551) xor estimated(555) xor estimated(559);
partial_sums(5)(402) <= estimated(291) xor estimated(295) xor estimated(299) xor estimated(303);
partial_sums(5)(403) <= estimated(803) xor estimated(807) xor estimated(811) xor estimated(815);
partial_sums(5)(404) <= estimated(163) xor estimated(167) xor estimated(171) xor estimated(175);
partial_sums(5)(405) <= estimated(675) xor estimated(679) xor estimated(683) xor estimated(687);
partial_sums(5)(406) <= estimated(419) xor estimated(423) xor estimated(427) xor estimated(431);
partial_sums(5)(407) <= estimated(931) xor estimated(935) xor estimated(939) xor estimated(943);
partial_sums(5)(408) <= estimated(99) xor estimated(103) xor estimated(107) xor estimated(111);
partial_sums(5)(409) <= estimated(611) xor estimated(615) xor estimated(619) xor estimated(623);
partial_sums(5)(410) <= estimated(355) xor estimated(359) xor estimated(363) xor estimated(367);
partial_sums(5)(411) <= estimated(867) xor estimated(871) xor estimated(875) xor estimated(879);
partial_sums(5)(412) <= estimated(227) xor estimated(231) xor estimated(235) xor estimated(239);
partial_sums(5)(413) <= estimated(739) xor estimated(743) xor estimated(747) xor estimated(751);
partial_sums(5)(414) <= estimated(483) xor estimated(487) xor estimated(491) xor estimated(495);
partial_sums(5)(415) <= estimated(995) xor estimated(999) xor estimated(1003) xor estimated(1007);
partial_sums(5)(416) <= estimated(11) xor estimated(15);
partial_sums(5)(417) <= estimated(523) xor estimated(527);
partial_sums(5)(418) <= estimated(267) xor estimated(271);
partial_sums(5)(419) <= estimated(779) xor estimated(783);
partial_sums(5)(420) <= estimated(139) xor estimated(143);
partial_sums(5)(421) <= estimated(651) xor estimated(655);
partial_sums(5)(422) <= estimated(395) xor estimated(399);
partial_sums(5)(423) <= estimated(907) xor estimated(911);
partial_sums(5)(424) <= estimated(75) xor estimated(79);
partial_sums(5)(425) <= estimated(587) xor estimated(591);
partial_sums(5)(426) <= estimated(331) xor estimated(335);
partial_sums(5)(427) <= estimated(843) xor estimated(847);
partial_sums(5)(428) <= estimated(203) xor estimated(207);
partial_sums(5)(429) <= estimated(715) xor estimated(719);
partial_sums(5)(430) <= estimated(459) xor estimated(463);
partial_sums(5)(431) <= estimated(971) xor estimated(975);
partial_sums(5)(432) <= estimated(43) xor estimated(47);
partial_sums(5)(433) <= estimated(555) xor estimated(559);
partial_sums(5)(434) <= estimated(299) xor estimated(303);
partial_sums(5)(435) <= estimated(811) xor estimated(815);
partial_sums(5)(436) <= estimated(171) xor estimated(175);
partial_sums(5)(437) <= estimated(683) xor estimated(687);
partial_sums(5)(438) <= estimated(427) xor estimated(431);
partial_sums(5)(439) <= estimated(939) xor estimated(943);
partial_sums(5)(440) <= estimated(107) xor estimated(111);
partial_sums(5)(441) <= estimated(619) xor estimated(623);
partial_sums(5)(442) <= estimated(363) xor estimated(367);
partial_sums(5)(443) <= estimated(875) xor estimated(879);
partial_sums(5)(444) <= estimated(235) xor estimated(239);
partial_sums(5)(445) <= estimated(747) xor estimated(751);
partial_sums(5)(446) <= estimated(491) xor estimated(495);
partial_sums(5)(447) <= estimated(1003) xor estimated(1007);
partial_sums(5)(448) <= estimated(7) xor estimated(15);
partial_sums(5)(449) <= estimated(519) xor estimated(527);
partial_sums(5)(450) <= estimated(263) xor estimated(271);
partial_sums(5)(451) <= estimated(775) xor estimated(783);
partial_sums(5)(452) <= estimated(135) xor estimated(143);
partial_sums(5)(453) <= estimated(647) xor estimated(655);
partial_sums(5)(454) <= estimated(391) xor estimated(399);
partial_sums(5)(455) <= estimated(903) xor estimated(911);
partial_sums(5)(456) <= estimated(71) xor estimated(79);
partial_sums(5)(457) <= estimated(583) xor estimated(591);
partial_sums(5)(458) <= estimated(327) xor estimated(335);
partial_sums(5)(459) <= estimated(839) xor estimated(847);
partial_sums(5)(460) <= estimated(199) xor estimated(207);
partial_sums(5)(461) <= estimated(711) xor estimated(719);
partial_sums(5)(462) <= estimated(455) xor estimated(463);
partial_sums(5)(463) <= estimated(967) xor estimated(975);
partial_sums(5)(464) <= estimated(39) xor estimated(47);
partial_sums(5)(465) <= estimated(551) xor estimated(559);
partial_sums(5)(466) <= estimated(295) xor estimated(303);
partial_sums(5)(467) <= estimated(807) xor estimated(815);
partial_sums(5)(468) <= estimated(167) xor estimated(175);
partial_sums(5)(469) <= estimated(679) xor estimated(687);
partial_sums(5)(470) <= estimated(423) xor estimated(431);
partial_sums(5)(471) <= estimated(935) xor estimated(943);
partial_sums(5)(472) <= estimated(103) xor estimated(111);
partial_sums(5)(473) <= estimated(615) xor estimated(623);
partial_sums(5)(474) <= estimated(359) xor estimated(367);
partial_sums(5)(475) <= estimated(871) xor estimated(879);
partial_sums(5)(476) <= estimated(231) xor estimated(239);
partial_sums(5)(477) <= estimated(743) xor estimated(751);
partial_sums(5)(478) <= estimated(487) xor estimated(495);
partial_sums(5)(479) <= estimated(999) xor estimated(1007);
partial_sums(5)(480) <= estimated(15);
partial_sums(5)(481) <= estimated(527);
partial_sums(5)(482) <= estimated(271);
partial_sums(5)(483) <= estimated(783);
partial_sums(5)(484) <= estimated(143);
partial_sums(5)(485) <= estimated(655);
partial_sums(5)(486) <= estimated(399);
partial_sums(5)(487) <= estimated(911);
partial_sums(5)(488) <= estimated(79);
partial_sums(5)(489) <= estimated(591);
partial_sums(5)(490) <= estimated(335);
partial_sums(5)(491) <= estimated(847);
partial_sums(5)(492) <= estimated(207);
partial_sums(5)(493) <= estimated(719);
partial_sums(5)(494) <= estimated(463);
partial_sums(5)(495) <= estimated(975);
partial_sums(5)(496) <= estimated(47);
partial_sums(5)(497) <= estimated(559);
partial_sums(5)(498) <= estimated(303);
partial_sums(5)(499) <= estimated(815);
partial_sums(5)(500) <= estimated(175);
partial_sums(5)(501) <= estimated(687);
partial_sums(5)(502) <= estimated(431);
partial_sums(5)(503) <= estimated(943);
partial_sums(5)(504) <= estimated(111);
partial_sums(5)(505) <= estimated(623);
partial_sums(5)(506) <= estimated(367);
partial_sums(5)(507) <= estimated(879);
partial_sums(5)(508) <= estimated(239);
partial_sums(5)(509) <= estimated(751);
partial_sums(5)(510) <= estimated(495);
partial_sums(5)(511) <= estimated(1007);
partial_sums(6)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(1) <= estimated(512) xor estimated(513) xor estimated(514) xor estimated(515) xor estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(2) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(3) <= estimated(768) xor estimated(769) xor estimated(770) xor estimated(771) xor estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(784) xor estimated(785) xor estimated(786) xor estimated(787) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(4) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(5) <= estimated(640) xor estimated(641) xor estimated(642) xor estimated(643) xor estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(6) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(7) <= estimated(896) xor estimated(897) xor estimated(898) xor estimated(899) xor estimated(900) xor estimated(901) xor estimated(902) xor estimated(903) xor estimated(904) xor estimated(905) xor estimated(906) xor estimated(907) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(912) xor estimated(913) xor estimated(914) xor estimated(915) xor estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(8) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(9) <= estimated(576) xor estimated(577) xor estimated(578) xor estimated(579) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(10) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(11) <= estimated(832) xor estimated(833) xor estimated(834) xor estimated(835) xor estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(848) xor estimated(849) xor estimated(850) xor estimated(851) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(12) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(13) <= estimated(704) xor estimated(705) xor estimated(706) xor estimated(707) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(14) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(15) <= estimated(960) xor estimated(961) xor estimated(962) xor estimated(963) xor estimated(964) xor estimated(965) xor estimated(966) xor estimated(967) xor estimated(968) xor estimated(969) xor estimated(970) xor estimated(971) xor estimated(972) xor estimated(973) xor estimated(974) xor estimated(975) xor estimated(976) xor estimated(977) xor estimated(978) xor estimated(979) xor estimated(980) xor estimated(981) xor estimated(982) xor estimated(983) xor estimated(984) xor estimated(985) xor estimated(986) xor estimated(987) xor estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(16) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(17) <= estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(18) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(19) <= estimated(784) xor estimated(785) xor estimated(786) xor estimated(787) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(20) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(21) <= estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(22) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(23) <= estimated(912) xor estimated(913) xor estimated(914) xor estimated(915) xor estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(24) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(25) <= estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(26) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(27) <= estimated(848) xor estimated(849) xor estimated(850) xor estimated(851) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(28) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(29) <= estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(30) <= estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(31) <= estimated(976) xor estimated(977) xor estimated(978) xor estimated(979) xor estimated(980) xor estimated(981) xor estimated(982) xor estimated(983) xor estimated(984) xor estimated(985) xor estimated(986) xor estimated(987) xor estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(32) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(33) <= estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(34) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(35) <= estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(36) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(37) <= estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(38) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(39) <= estimated(904) xor estimated(905) xor estimated(906) xor estimated(907) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(40) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(41) <= estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(42) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(43) <= estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(44) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(45) <= estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(46) <= estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(47) <= estimated(968) xor estimated(969) xor estimated(970) xor estimated(971) xor estimated(972) xor estimated(973) xor estimated(974) xor estimated(975) xor estimated(984) xor estimated(985) xor estimated(986) xor estimated(987) xor estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(48) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(49) <= estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(50) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(51) <= estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(52) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(53) <= estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(54) <= estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(55) <= estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(56) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(57) <= estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(58) <= estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(59) <= estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(60) <= estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(61) <= estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(62) <= estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(63) <= estimated(984) xor estimated(985) xor estimated(986) xor estimated(987) xor estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(64) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(65) <= estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(66) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(67) <= estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(68) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(69) <= estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(70) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(71) <= estimated(900) xor estimated(901) xor estimated(902) xor estimated(903) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(72) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(73) <= estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(74) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(75) <= estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(76) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(77) <= estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(78) <= estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(79) <= estimated(964) xor estimated(965) xor estimated(966) xor estimated(967) xor estimated(972) xor estimated(973) xor estimated(974) xor estimated(975) xor estimated(980) xor estimated(981) xor estimated(982) xor estimated(983) xor estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(80) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(81) <= estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(82) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(83) <= estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(84) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(85) <= estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(86) <= estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(87) <= estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(88) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(89) <= estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(90) <= estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(91) <= estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(92) <= estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(93) <= estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(94) <= estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(95) <= estimated(980) xor estimated(981) xor estimated(982) xor estimated(983) xor estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(96) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(97) <= estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(98) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(99) <= estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(100) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(101) <= estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(102) <= estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(103) <= estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(104) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(105) <= estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(106) <= estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(107) <= estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(108) <= estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(109) <= estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(110) <= estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(111) <= estimated(972) xor estimated(973) xor estimated(974) xor estimated(975) xor estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(112) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31);
partial_sums(6)(113) <= estimated(540) xor estimated(541) xor estimated(542) xor estimated(543);
partial_sums(6)(114) <= estimated(284) xor estimated(285) xor estimated(286) xor estimated(287);
partial_sums(6)(115) <= estimated(796) xor estimated(797) xor estimated(798) xor estimated(799);
partial_sums(6)(116) <= estimated(156) xor estimated(157) xor estimated(158) xor estimated(159);
partial_sums(6)(117) <= estimated(668) xor estimated(669) xor estimated(670) xor estimated(671);
partial_sums(6)(118) <= estimated(412) xor estimated(413) xor estimated(414) xor estimated(415);
partial_sums(6)(119) <= estimated(924) xor estimated(925) xor estimated(926) xor estimated(927);
partial_sums(6)(120) <= estimated(92) xor estimated(93) xor estimated(94) xor estimated(95);
partial_sums(6)(121) <= estimated(604) xor estimated(605) xor estimated(606) xor estimated(607);
partial_sums(6)(122) <= estimated(348) xor estimated(349) xor estimated(350) xor estimated(351);
partial_sums(6)(123) <= estimated(860) xor estimated(861) xor estimated(862) xor estimated(863);
partial_sums(6)(124) <= estimated(220) xor estimated(221) xor estimated(222) xor estimated(223);
partial_sums(6)(125) <= estimated(732) xor estimated(733) xor estimated(734) xor estimated(735);
partial_sums(6)(126) <= estimated(476) xor estimated(477) xor estimated(478) xor estimated(479);
partial_sums(6)(127) <= estimated(988) xor estimated(989) xor estimated(990) xor estimated(991);
partial_sums(6)(128) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(129) <= estimated(514) xor estimated(515) xor estimated(518) xor estimated(519) xor estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543);
partial_sums(6)(130) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(131) <= estimated(770) xor estimated(771) xor estimated(774) xor estimated(775) xor estimated(778) xor estimated(779) xor estimated(782) xor estimated(783) xor estimated(786) xor estimated(787) xor estimated(790) xor estimated(791) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799);
partial_sums(6)(132) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(133) <= estimated(642) xor estimated(643) xor estimated(646) xor estimated(647) xor estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671);
partial_sums(6)(134) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(135) <= estimated(898) xor estimated(899) xor estimated(902) xor estimated(903) xor estimated(906) xor estimated(907) xor estimated(910) xor estimated(911) xor estimated(914) xor estimated(915) xor estimated(918) xor estimated(919) xor estimated(922) xor estimated(923) xor estimated(926) xor estimated(927);
partial_sums(6)(136) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(137) <= estimated(578) xor estimated(579) xor estimated(582) xor estimated(583) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607);
partial_sums(6)(138) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(139) <= estimated(834) xor estimated(835) xor estimated(838) xor estimated(839) xor estimated(842) xor estimated(843) xor estimated(846) xor estimated(847) xor estimated(850) xor estimated(851) xor estimated(854) xor estimated(855) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863);
partial_sums(6)(140) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(141) <= estimated(706) xor estimated(707) xor estimated(710) xor estimated(711) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735);
partial_sums(6)(142) <= estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(143) <= estimated(962) xor estimated(963) xor estimated(966) xor estimated(967) xor estimated(970) xor estimated(971) xor estimated(974) xor estimated(975) xor estimated(978) xor estimated(979) xor estimated(982) xor estimated(983) xor estimated(986) xor estimated(987) xor estimated(990) xor estimated(991);
partial_sums(6)(144) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(145) <= estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543);
partial_sums(6)(146) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(147) <= estimated(786) xor estimated(787) xor estimated(790) xor estimated(791) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799);
partial_sums(6)(148) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(149) <= estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671);
partial_sums(6)(150) <= estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(151) <= estimated(914) xor estimated(915) xor estimated(918) xor estimated(919) xor estimated(922) xor estimated(923) xor estimated(926) xor estimated(927);
partial_sums(6)(152) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(153) <= estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607);
partial_sums(6)(154) <= estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(155) <= estimated(850) xor estimated(851) xor estimated(854) xor estimated(855) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863);
partial_sums(6)(156) <= estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(157) <= estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735);
partial_sums(6)(158) <= estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(159) <= estimated(978) xor estimated(979) xor estimated(982) xor estimated(983) xor estimated(986) xor estimated(987) xor estimated(990) xor estimated(991);
partial_sums(6)(160) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(161) <= estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543);
partial_sums(6)(162) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(163) <= estimated(778) xor estimated(779) xor estimated(782) xor estimated(783) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799);
partial_sums(6)(164) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(165) <= estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671);
partial_sums(6)(166) <= estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(167) <= estimated(906) xor estimated(907) xor estimated(910) xor estimated(911) xor estimated(922) xor estimated(923) xor estimated(926) xor estimated(927);
partial_sums(6)(168) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(169) <= estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607);
partial_sums(6)(170) <= estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(171) <= estimated(842) xor estimated(843) xor estimated(846) xor estimated(847) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863);
partial_sums(6)(172) <= estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(173) <= estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735);
partial_sums(6)(174) <= estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(175) <= estimated(970) xor estimated(971) xor estimated(974) xor estimated(975) xor estimated(986) xor estimated(987) xor estimated(990) xor estimated(991);
partial_sums(6)(176) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31);
partial_sums(6)(177) <= estimated(538) xor estimated(539) xor estimated(542) xor estimated(543);
partial_sums(6)(178) <= estimated(282) xor estimated(283) xor estimated(286) xor estimated(287);
partial_sums(6)(179) <= estimated(794) xor estimated(795) xor estimated(798) xor estimated(799);
partial_sums(6)(180) <= estimated(154) xor estimated(155) xor estimated(158) xor estimated(159);
partial_sums(6)(181) <= estimated(666) xor estimated(667) xor estimated(670) xor estimated(671);
partial_sums(6)(182) <= estimated(410) xor estimated(411) xor estimated(414) xor estimated(415);
partial_sums(6)(183) <= estimated(922) xor estimated(923) xor estimated(926) xor estimated(927);
partial_sums(6)(184) <= estimated(90) xor estimated(91) xor estimated(94) xor estimated(95);
partial_sums(6)(185) <= estimated(602) xor estimated(603) xor estimated(606) xor estimated(607);
partial_sums(6)(186) <= estimated(346) xor estimated(347) xor estimated(350) xor estimated(351);
partial_sums(6)(187) <= estimated(858) xor estimated(859) xor estimated(862) xor estimated(863);
partial_sums(6)(188) <= estimated(218) xor estimated(219) xor estimated(222) xor estimated(223);
partial_sums(6)(189) <= estimated(730) xor estimated(731) xor estimated(734) xor estimated(735);
partial_sums(6)(190) <= estimated(474) xor estimated(475) xor estimated(478) xor estimated(479);
partial_sums(6)(191) <= estimated(986) xor estimated(987) xor estimated(990) xor estimated(991);
partial_sums(6)(192) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31);
partial_sums(6)(193) <= estimated(518) xor estimated(519) xor estimated(526) xor estimated(527) xor estimated(534) xor estimated(535) xor estimated(542) xor estimated(543);
partial_sums(6)(194) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287);
partial_sums(6)(195) <= estimated(774) xor estimated(775) xor estimated(782) xor estimated(783) xor estimated(790) xor estimated(791) xor estimated(798) xor estimated(799);
partial_sums(6)(196) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159);
partial_sums(6)(197) <= estimated(646) xor estimated(647) xor estimated(654) xor estimated(655) xor estimated(662) xor estimated(663) xor estimated(670) xor estimated(671);
partial_sums(6)(198) <= estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415);
partial_sums(6)(199) <= estimated(902) xor estimated(903) xor estimated(910) xor estimated(911) xor estimated(918) xor estimated(919) xor estimated(926) xor estimated(927);
partial_sums(6)(200) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95);
partial_sums(6)(201) <= estimated(582) xor estimated(583) xor estimated(590) xor estimated(591) xor estimated(598) xor estimated(599) xor estimated(606) xor estimated(607);
partial_sums(6)(202) <= estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351);
partial_sums(6)(203) <= estimated(838) xor estimated(839) xor estimated(846) xor estimated(847) xor estimated(854) xor estimated(855) xor estimated(862) xor estimated(863);
partial_sums(6)(204) <= estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223);
partial_sums(6)(205) <= estimated(710) xor estimated(711) xor estimated(718) xor estimated(719) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735);
partial_sums(6)(206) <= estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479);
partial_sums(6)(207) <= estimated(966) xor estimated(967) xor estimated(974) xor estimated(975) xor estimated(982) xor estimated(983) xor estimated(990) xor estimated(991);
partial_sums(6)(208) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31);
partial_sums(6)(209) <= estimated(534) xor estimated(535) xor estimated(542) xor estimated(543);
partial_sums(6)(210) <= estimated(278) xor estimated(279) xor estimated(286) xor estimated(287);
partial_sums(6)(211) <= estimated(790) xor estimated(791) xor estimated(798) xor estimated(799);
partial_sums(6)(212) <= estimated(150) xor estimated(151) xor estimated(158) xor estimated(159);
partial_sums(6)(213) <= estimated(662) xor estimated(663) xor estimated(670) xor estimated(671);
partial_sums(6)(214) <= estimated(406) xor estimated(407) xor estimated(414) xor estimated(415);
partial_sums(6)(215) <= estimated(918) xor estimated(919) xor estimated(926) xor estimated(927);
partial_sums(6)(216) <= estimated(86) xor estimated(87) xor estimated(94) xor estimated(95);
partial_sums(6)(217) <= estimated(598) xor estimated(599) xor estimated(606) xor estimated(607);
partial_sums(6)(218) <= estimated(342) xor estimated(343) xor estimated(350) xor estimated(351);
partial_sums(6)(219) <= estimated(854) xor estimated(855) xor estimated(862) xor estimated(863);
partial_sums(6)(220) <= estimated(214) xor estimated(215) xor estimated(222) xor estimated(223);
partial_sums(6)(221) <= estimated(726) xor estimated(727) xor estimated(734) xor estimated(735);
partial_sums(6)(222) <= estimated(470) xor estimated(471) xor estimated(478) xor estimated(479);
partial_sums(6)(223) <= estimated(982) xor estimated(983) xor estimated(990) xor estimated(991);
partial_sums(6)(224) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31);
partial_sums(6)(225) <= estimated(526) xor estimated(527) xor estimated(542) xor estimated(543);
partial_sums(6)(226) <= estimated(270) xor estimated(271) xor estimated(286) xor estimated(287);
partial_sums(6)(227) <= estimated(782) xor estimated(783) xor estimated(798) xor estimated(799);
partial_sums(6)(228) <= estimated(142) xor estimated(143) xor estimated(158) xor estimated(159);
partial_sums(6)(229) <= estimated(654) xor estimated(655) xor estimated(670) xor estimated(671);
partial_sums(6)(230) <= estimated(398) xor estimated(399) xor estimated(414) xor estimated(415);
partial_sums(6)(231) <= estimated(910) xor estimated(911) xor estimated(926) xor estimated(927);
partial_sums(6)(232) <= estimated(78) xor estimated(79) xor estimated(94) xor estimated(95);
partial_sums(6)(233) <= estimated(590) xor estimated(591) xor estimated(606) xor estimated(607);
partial_sums(6)(234) <= estimated(334) xor estimated(335) xor estimated(350) xor estimated(351);
partial_sums(6)(235) <= estimated(846) xor estimated(847) xor estimated(862) xor estimated(863);
partial_sums(6)(236) <= estimated(206) xor estimated(207) xor estimated(222) xor estimated(223);
partial_sums(6)(237) <= estimated(718) xor estimated(719) xor estimated(734) xor estimated(735);
partial_sums(6)(238) <= estimated(462) xor estimated(463) xor estimated(478) xor estimated(479);
partial_sums(6)(239) <= estimated(974) xor estimated(975) xor estimated(990) xor estimated(991);
partial_sums(6)(240) <= estimated(30) xor estimated(31);
partial_sums(6)(241) <= estimated(542) xor estimated(543);
partial_sums(6)(242) <= estimated(286) xor estimated(287);
partial_sums(6)(243) <= estimated(798) xor estimated(799);
partial_sums(6)(244) <= estimated(158) xor estimated(159);
partial_sums(6)(245) <= estimated(670) xor estimated(671);
partial_sums(6)(246) <= estimated(414) xor estimated(415);
partial_sums(6)(247) <= estimated(926) xor estimated(927);
partial_sums(6)(248) <= estimated(94) xor estimated(95);
partial_sums(6)(249) <= estimated(606) xor estimated(607);
partial_sums(6)(250) <= estimated(350) xor estimated(351);
partial_sums(6)(251) <= estimated(862) xor estimated(863);
partial_sums(6)(252) <= estimated(222) xor estimated(223);
partial_sums(6)(253) <= estimated(734) xor estimated(735);
partial_sums(6)(254) <= estimated(478) xor estimated(479);
partial_sums(6)(255) <= estimated(990) xor estimated(991);
partial_sums(6)(256) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(257) <= estimated(513) xor estimated(515) xor estimated(517) xor estimated(519) xor estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543);
partial_sums(6)(258) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(259) <= estimated(769) xor estimated(771) xor estimated(773) xor estimated(775) xor estimated(777) xor estimated(779) xor estimated(781) xor estimated(783) xor estimated(785) xor estimated(787) xor estimated(789) xor estimated(791) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799);
partial_sums(6)(260) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(261) <= estimated(641) xor estimated(643) xor estimated(645) xor estimated(647) xor estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671);
partial_sums(6)(262) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(263) <= estimated(897) xor estimated(899) xor estimated(901) xor estimated(903) xor estimated(905) xor estimated(907) xor estimated(909) xor estimated(911) xor estimated(913) xor estimated(915) xor estimated(917) xor estimated(919) xor estimated(921) xor estimated(923) xor estimated(925) xor estimated(927);
partial_sums(6)(264) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(265) <= estimated(577) xor estimated(579) xor estimated(581) xor estimated(583) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607);
partial_sums(6)(266) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(267) <= estimated(833) xor estimated(835) xor estimated(837) xor estimated(839) xor estimated(841) xor estimated(843) xor estimated(845) xor estimated(847) xor estimated(849) xor estimated(851) xor estimated(853) xor estimated(855) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863);
partial_sums(6)(268) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(269) <= estimated(705) xor estimated(707) xor estimated(709) xor estimated(711) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735);
partial_sums(6)(270) <= estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(271) <= estimated(961) xor estimated(963) xor estimated(965) xor estimated(967) xor estimated(969) xor estimated(971) xor estimated(973) xor estimated(975) xor estimated(977) xor estimated(979) xor estimated(981) xor estimated(983) xor estimated(985) xor estimated(987) xor estimated(989) xor estimated(991);
partial_sums(6)(272) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(273) <= estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543);
partial_sums(6)(274) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(275) <= estimated(785) xor estimated(787) xor estimated(789) xor estimated(791) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799);
partial_sums(6)(276) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(277) <= estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671);
partial_sums(6)(278) <= estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(279) <= estimated(913) xor estimated(915) xor estimated(917) xor estimated(919) xor estimated(921) xor estimated(923) xor estimated(925) xor estimated(927);
partial_sums(6)(280) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(281) <= estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607);
partial_sums(6)(282) <= estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(283) <= estimated(849) xor estimated(851) xor estimated(853) xor estimated(855) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863);
partial_sums(6)(284) <= estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(285) <= estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735);
partial_sums(6)(286) <= estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(287) <= estimated(977) xor estimated(979) xor estimated(981) xor estimated(983) xor estimated(985) xor estimated(987) xor estimated(989) xor estimated(991);
partial_sums(6)(288) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(289) <= estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543);
partial_sums(6)(290) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(291) <= estimated(777) xor estimated(779) xor estimated(781) xor estimated(783) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799);
partial_sums(6)(292) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(293) <= estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671);
partial_sums(6)(294) <= estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(295) <= estimated(905) xor estimated(907) xor estimated(909) xor estimated(911) xor estimated(921) xor estimated(923) xor estimated(925) xor estimated(927);
partial_sums(6)(296) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(297) <= estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607);
partial_sums(6)(298) <= estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(299) <= estimated(841) xor estimated(843) xor estimated(845) xor estimated(847) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863);
partial_sums(6)(300) <= estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(301) <= estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735);
partial_sums(6)(302) <= estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(303) <= estimated(969) xor estimated(971) xor estimated(973) xor estimated(975) xor estimated(985) xor estimated(987) xor estimated(989) xor estimated(991);
partial_sums(6)(304) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31);
partial_sums(6)(305) <= estimated(537) xor estimated(539) xor estimated(541) xor estimated(543);
partial_sums(6)(306) <= estimated(281) xor estimated(283) xor estimated(285) xor estimated(287);
partial_sums(6)(307) <= estimated(793) xor estimated(795) xor estimated(797) xor estimated(799);
partial_sums(6)(308) <= estimated(153) xor estimated(155) xor estimated(157) xor estimated(159);
partial_sums(6)(309) <= estimated(665) xor estimated(667) xor estimated(669) xor estimated(671);
partial_sums(6)(310) <= estimated(409) xor estimated(411) xor estimated(413) xor estimated(415);
partial_sums(6)(311) <= estimated(921) xor estimated(923) xor estimated(925) xor estimated(927);
partial_sums(6)(312) <= estimated(89) xor estimated(91) xor estimated(93) xor estimated(95);
partial_sums(6)(313) <= estimated(601) xor estimated(603) xor estimated(605) xor estimated(607);
partial_sums(6)(314) <= estimated(345) xor estimated(347) xor estimated(349) xor estimated(351);
partial_sums(6)(315) <= estimated(857) xor estimated(859) xor estimated(861) xor estimated(863);
partial_sums(6)(316) <= estimated(217) xor estimated(219) xor estimated(221) xor estimated(223);
partial_sums(6)(317) <= estimated(729) xor estimated(731) xor estimated(733) xor estimated(735);
partial_sums(6)(318) <= estimated(473) xor estimated(475) xor estimated(477) xor estimated(479);
partial_sums(6)(319) <= estimated(985) xor estimated(987) xor estimated(989) xor estimated(991);
partial_sums(6)(320) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31);
partial_sums(6)(321) <= estimated(517) xor estimated(519) xor estimated(525) xor estimated(527) xor estimated(533) xor estimated(535) xor estimated(541) xor estimated(543);
partial_sums(6)(322) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287);
partial_sums(6)(323) <= estimated(773) xor estimated(775) xor estimated(781) xor estimated(783) xor estimated(789) xor estimated(791) xor estimated(797) xor estimated(799);
partial_sums(6)(324) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159);
partial_sums(6)(325) <= estimated(645) xor estimated(647) xor estimated(653) xor estimated(655) xor estimated(661) xor estimated(663) xor estimated(669) xor estimated(671);
partial_sums(6)(326) <= estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415);
partial_sums(6)(327) <= estimated(901) xor estimated(903) xor estimated(909) xor estimated(911) xor estimated(917) xor estimated(919) xor estimated(925) xor estimated(927);
partial_sums(6)(328) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95);
partial_sums(6)(329) <= estimated(581) xor estimated(583) xor estimated(589) xor estimated(591) xor estimated(597) xor estimated(599) xor estimated(605) xor estimated(607);
partial_sums(6)(330) <= estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351);
partial_sums(6)(331) <= estimated(837) xor estimated(839) xor estimated(845) xor estimated(847) xor estimated(853) xor estimated(855) xor estimated(861) xor estimated(863);
partial_sums(6)(332) <= estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223);
partial_sums(6)(333) <= estimated(709) xor estimated(711) xor estimated(717) xor estimated(719) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735);
partial_sums(6)(334) <= estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479);
partial_sums(6)(335) <= estimated(965) xor estimated(967) xor estimated(973) xor estimated(975) xor estimated(981) xor estimated(983) xor estimated(989) xor estimated(991);
partial_sums(6)(336) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31);
partial_sums(6)(337) <= estimated(533) xor estimated(535) xor estimated(541) xor estimated(543);
partial_sums(6)(338) <= estimated(277) xor estimated(279) xor estimated(285) xor estimated(287);
partial_sums(6)(339) <= estimated(789) xor estimated(791) xor estimated(797) xor estimated(799);
partial_sums(6)(340) <= estimated(149) xor estimated(151) xor estimated(157) xor estimated(159);
partial_sums(6)(341) <= estimated(661) xor estimated(663) xor estimated(669) xor estimated(671);
partial_sums(6)(342) <= estimated(405) xor estimated(407) xor estimated(413) xor estimated(415);
partial_sums(6)(343) <= estimated(917) xor estimated(919) xor estimated(925) xor estimated(927);
partial_sums(6)(344) <= estimated(85) xor estimated(87) xor estimated(93) xor estimated(95);
partial_sums(6)(345) <= estimated(597) xor estimated(599) xor estimated(605) xor estimated(607);
partial_sums(6)(346) <= estimated(341) xor estimated(343) xor estimated(349) xor estimated(351);
partial_sums(6)(347) <= estimated(853) xor estimated(855) xor estimated(861) xor estimated(863);
partial_sums(6)(348) <= estimated(213) xor estimated(215) xor estimated(221) xor estimated(223);
partial_sums(6)(349) <= estimated(725) xor estimated(727) xor estimated(733) xor estimated(735);
partial_sums(6)(350) <= estimated(469) xor estimated(471) xor estimated(477) xor estimated(479);
partial_sums(6)(351) <= estimated(981) xor estimated(983) xor estimated(989) xor estimated(991);
partial_sums(6)(352) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31);
partial_sums(6)(353) <= estimated(525) xor estimated(527) xor estimated(541) xor estimated(543);
partial_sums(6)(354) <= estimated(269) xor estimated(271) xor estimated(285) xor estimated(287);
partial_sums(6)(355) <= estimated(781) xor estimated(783) xor estimated(797) xor estimated(799);
partial_sums(6)(356) <= estimated(141) xor estimated(143) xor estimated(157) xor estimated(159);
partial_sums(6)(357) <= estimated(653) xor estimated(655) xor estimated(669) xor estimated(671);
partial_sums(6)(358) <= estimated(397) xor estimated(399) xor estimated(413) xor estimated(415);
partial_sums(6)(359) <= estimated(909) xor estimated(911) xor estimated(925) xor estimated(927);
partial_sums(6)(360) <= estimated(77) xor estimated(79) xor estimated(93) xor estimated(95);
partial_sums(6)(361) <= estimated(589) xor estimated(591) xor estimated(605) xor estimated(607);
partial_sums(6)(362) <= estimated(333) xor estimated(335) xor estimated(349) xor estimated(351);
partial_sums(6)(363) <= estimated(845) xor estimated(847) xor estimated(861) xor estimated(863);
partial_sums(6)(364) <= estimated(205) xor estimated(207) xor estimated(221) xor estimated(223);
partial_sums(6)(365) <= estimated(717) xor estimated(719) xor estimated(733) xor estimated(735);
partial_sums(6)(366) <= estimated(461) xor estimated(463) xor estimated(477) xor estimated(479);
partial_sums(6)(367) <= estimated(973) xor estimated(975) xor estimated(989) xor estimated(991);
partial_sums(6)(368) <= estimated(29) xor estimated(31);
partial_sums(6)(369) <= estimated(541) xor estimated(543);
partial_sums(6)(370) <= estimated(285) xor estimated(287);
partial_sums(6)(371) <= estimated(797) xor estimated(799);
partial_sums(6)(372) <= estimated(157) xor estimated(159);
partial_sums(6)(373) <= estimated(669) xor estimated(671);
partial_sums(6)(374) <= estimated(413) xor estimated(415);
partial_sums(6)(375) <= estimated(925) xor estimated(927);
partial_sums(6)(376) <= estimated(93) xor estimated(95);
partial_sums(6)(377) <= estimated(605) xor estimated(607);
partial_sums(6)(378) <= estimated(349) xor estimated(351);
partial_sums(6)(379) <= estimated(861) xor estimated(863);
partial_sums(6)(380) <= estimated(221) xor estimated(223);
partial_sums(6)(381) <= estimated(733) xor estimated(735);
partial_sums(6)(382) <= estimated(477) xor estimated(479);
partial_sums(6)(383) <= estimated(989) xor estimated(991);
partial_sums(6)(384) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31);
partial_sums(6)(385) <= estimated(515) xor estimated(519) xor estimated(523) xor estimated(527) xor estimated(531) xor estimated(535) xor estimated(539) xor estimated(543);
partial_sums(6)(386) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287);
partial_sums(6)(387) <= estimated(771) xor estimated(775) xor estimated(779) xor estimated(783) xor estimated(787) xor estimated(791) xor estimated(795) xor estimated(799);
partial_sums(6)(388) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159);
partial_sums(6)(389) <= estimated(643) xor estimated(647) xor estimated(651) xor estimated(655) xor estimated(659) xor estimated(663) xor estimated(667) xor estimated(671);
partial_sums(6)(390) <= estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415);
partial_sums(6)(391) <= estimated(899) xor estimated(903) xor estimated(907) xor estimated(911) xor estimated(915) xor estimated(919) xor estimated(923) xor estimated(927);
partial_sums(6)(392) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95);
partial_sums(6)(393) <= estimated(579) xor estimated(583) xor estimated(587) xor estimated(591) xor estimated(595) xor estimated(599) xor estimated(603) xor estimated(607);
partial_sums(6)(394) <= estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351);
partial_sums(6)(395) <= estimated(835) xor estimated(839) xor estimated(843) xor estimated(847) xor estimated(851) xor estimated(855) xor estimated(859) xor estimated(863);
partial_sums(6)(396) <= estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223);
partial_sums(6)(397) <= estimated(707) xor estimated(711) xor estimated(715) xor estimated(719) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735);
partial_sums(6)(398) <= estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479);
partial_sums(6)(399) <= estimated(963) xor estimated(967) xor estimated(971) xor estimated(975) xor estimated(979) xor estimated(983) xor estimated(987) xor estimated(991);
partial_sums(6)(400) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31);
partial_sums(6)(401) <= estimated(531) xor estimated(535) xor estimated(539) xor estimated(543);
partial_sums(6)(402) <= estimated(275) xor estimated(279) xor estimated(283) xor estimated(287);
partial_sums(6)(403) <= estimated(787) xor estimated(791) xor estimated(795) xor estimated(799);
partial_sums(6)(404) <= estimated(147) xor estimated(151) xor estimated(155) xor estimated(159);
partial_sums(6)(405) <= estimated(659) xor estimated(663) xor estimated(667) xor estimated(671);
partial_sums(6)(406) <= estimated(403) xor estimated(407) xor estimated(411) xor estimated(415);
partial_sums(6)(407) <= estimated(915) xor estimated(919) xor estimated(923) xor estimated(927);
partial_sums(6)(408) <= estimated(83) xor estimated(87) xor estimated(91) xor estimated(95);
partial_sums(6)(409) <= estimated(595) xor estimated(599) xor estimated(603) xor estimated(607);
partial_sums(6)(410) <= estimated(339) xor estimated(343) xor estimated(347) xor estimated(351);
partial_sums(6)(411) <= estimated(851) xor estimated(855) xor estimated(859) xor estimated(863);
partial_sums(6)(412) <= estimated(211) xor estimated(215) xor estimated(219) xor estimated(223);
partial_sums(6)(413) <= estimated(723) xor estimated(727) xor estimated(731) xor estimated(735);
partial_sums(6)(414) <= estimated(467) xor estimated(471) xor estimated(475) xor estimated(479);
partial_sums(6)(415) <= estimated(979) xor estimated(983) xor estimated(987) xor estimated(991);
partial_sums(6)(416) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31);
partial_sums(6)(417) <= estimated(523) xor estimated(527) xor estimated(539) xor estimated(543);
partial_sums(6)(418) <= estimated(267) xor estimated(271) xor estimated(283) xor estimated(287);
partial_sums(6)(419) <= estimated(779) xor estimated(783) xor estimated(795) xor estimated(799);
partial_sums(6)(420) <= estimated(139) xor estimated(143) xor estimated(155) xor estimated(159);
partial_sums(6)(421) <= estimated(651) xor estimated(655) xor estimated(667) xor estimated(671);
partial_sums(6)(422) <= estimated(395) xor estimated(399) xor estimated(411) xor estimated(415);
partial_sums(6)(423) <= estimated(907) xor estimated(911) xor estimated(923) xor estimated(927);
partial_sums(6)(424) <= estimated(75) xor estimated(79) xor estimated(91) xor estimated(95);
partial_sums(6)(425) <= estimated(587) xor estimated(591) xor estimated(603) xor estimated(607);
partial_sums(6)(426) <= estimated(331) xor estimated(335) xor estimated(347) xor estimated(351);
partial_sums(6)(427) <= estimated(843) xor estimated(847) xor estimated(859) xor estimated(863);
partial_sums(6)(428) <= estimated(203) xor estimated(207) xor estimated(219) xor estimated(223);
partial_sums(6)(429) <= estimated(715) xor estimated(719) xor estimated(731) xor estimated(735);
partial_sums(6)(430) <= estimated(459) xor estimated(463) xor estimated(475) xor estimated(479);
partial_sums(6)(431) <= estimated(971) xor estimated(975) xor estimated(987) xor estimated(991);
partial_sums(6)(432) <= estimated(27) xor estimated(31);
partial_sums(6)(433) <= estimated(539) xor estimated(543);
partial_sums(6)(434) <= estimated(283) xor estimated(287);
partial_sums(6)(435) <= estimated(795) xor estimated(799);
partial_sums(6)(436) <= estimated(155) xor estimated(159);
partial_sums(6)(437) <= estimated(667) xor estimated(671);
partial_sums(6)(438) <= estimated(411) xor estimated(415);
partial_sums(6)(439) <= estimated(923) xor estimated(927);
partial_sums(6)(440) <= estimated(91) xor estimated(95);
partial_sums(6)(441) <= estimated(603) xor estimated(607);
partial_sums(6)(442) <= estimated(347) xor estimated(351);
partial_sums(6)(443) <= estimated(859) xor estimated(863);
partial_sums(6)(444) <= estimated(219) xor estimated(223);
partial_sums(6)(445) <= estimated(731) xor estimated(735);
partial_sums(6)(446) <= estimated(475) xor estimated(479);
partial_sums(6)(447) <= estimated(987) xor estimated(991);
partial_sums(6)(448) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31);
partial_sums(6)(449) <= estimated(519) xor estimated(527) xor estimated(535) xor estimated(543);
partial_sums(6)(450) <= estimated(263) xor estimated(271) xor estimated(279) xor estimated(287);
partial_sums(6)(451) <= estimated(775) xor estimated(783) xor estimated(791) xor estimated(799);
partial_sums(6)(452) <= estimated(135) xor estimated(143) xor estimated(151) xor estimated(159);
partial_sums(6)(453) <= estimated(647) xor estimated(655) xor estimated(663) xor estimated(671);
partial_sums(6)(454) <= estimated(391) xor estimated(399) xor estimated(407) xor estimated(415);
partial_sums(6)(455) <= estimated(903) xor estimated(911) xor estimated(919) xor estimated(927);
partial_sums(6)(456) <= estimated(71) xor estimated(79) xor estimated(87) xor estimated(95);
partial_sums(6)(457) <= estimated(583) xor estimated(591) xor estimated(599) xor estimated(607);
partial_sums(6)(458) <= estimated(327) xor estimated(335) xor estimated(343) xor estimated(351);
partial_sums(6)(459) <= estimated(839) xor estimated(847) xor estimated(855) xor estimated(863);
partial_sums(6)(460) <= estimated(199) xor estimated(207) xor estimated(215) xor estimated(223);
partial_sums(6)(461) <= estimated(711) xor estimated(719) xor estimated(727) xor estimated(735);
partial_sums(6)(462) <= estimated(455) xor estimated(463) xor estimated(471) xor estimated(479);
partial_sums(6)(463) <= estimated(967) xor estimated(975) xor estimated(983) xor estimated(991);
partial_sums(6)(464) <= estimated(23) xor estimated(31);
partial_sums(6)(465) <= estimated(535) xor estimated(543);
partial_sums(6)(466) <= estimated(279) xor estimated(287);
partial_sums(6)(467) <= estimated(791) xor estimated(799);
partial_sums(6)(468) <= estimated(151) xor estimated(159);
partial_sums(6)(469) <= estimated(663) xor estimated(671);
partial_sums(6)(470) <= estimated(407) xor estimated(415);
partial_sums(6)(471) <= estimated(919) xor estimated(927);
partial_sums(6)(472) <= estimated(87) xor estimated(95);
partial_sums(6)(473) <= estimated(599) xor estimated(607);
partial_sums(6)(474) <= estimated(343) xor estimated(351);
partial_sums(6)(475) <= estimated(855) xor estimated(863);
partial_sums(6)(476) <= estimated(215) xor estimated(223);
partial_sums(6)(477) <= estimated(727) xor estimated(735);
partial_sums(6)(478) <= estimated(471) xor estimated(479);
partial_sums(6)(479) <= estimated(983) xor estimated(991);
partial_sums(6)(480) <= estimated(15) xor estimated(31);
partial_sums(6)(481) <= estimated(527) xor estimated(543);
partial_sums(6)(482) <= estimated(271) xor estimated(287);
partial_sums(6)(483) <= estimated(783) xor estimated(799);
partial_sums(6)(484) <= estimated(143) xor estimated(159);
partial_sums(6)(485) <= estimated(655) xor estimated(671);
partial_sums(6)(486) <= estimated(399) xor estimated(415);
partial_sums(6)(487) <= estimated(911) xor estimated(927);
partial_sums(6)(488) <= estimated(79) xor estimated(95);
partial_sums(6)(489) <= estimated(591) xor estimated(607);
partial_sums(6)(490) <= estimated(335) xor estimated(351);
partial_sums(6)(491) <= estimated(847) xor estimated(863);
partial_sums(6)(492) <= estimated(207) xor estimated(223);
partial_sums(6)(493) <= estimated(719) xor estimated(735);
partial_sums(6)(494) <= estimated(463) xor estimated(479);
partial_sums(6)(495) <= estimated(975) xor estimated(991);
partial_sums(6)(496) <= estimated(31);
partial_sums(6)(497) <= estimated(543);
partial_sums(6)(498) <= estimated(287);
partial_sums(6)(499) <= estimated(799);
partial_sums(6)(500) <= estimated(159);
partial_sums(6)(501) <= estimated(671);
partial_sums(6)(502) <= estimated(415);
partial_sums(6)(503) <= estimated(927);
partial_sums(6)(504) <= estimated(95);
partial_sums(6)(505) <= estimated(607);
partial_sums(6)(506) <= estimated(351);
partial_sums(6)(507) <= estimated(863);
partial_sums(6)(508) <= estimated(223);
partial_sums(6)(509) <= estimated(735);
partial_sums(6)(510) <= estimated(479);
partial_sums(6)(511) <= estimated(991);
partial_sums(7)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(1) <= estimated(512) xor estimated(513) xor estimated(514) xor estimated(515) xor estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(2) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(3) <= estimated(768) xor estimated(769) xor estimated(770) xor estimated(771) xor estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(784) xor estimated(785) xor estimated(786) xor estimated(787) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(800) xor estimated(801) xor estimated(802) xor estimated(803) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(4) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(5) <= estimated(640) xor estimated(641) xor estimated(642) xor estimated(643) xor estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(6) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(7) <= estimated(896) xor estimated(897) xor estimated(898) xor estimated(899) xor estimated(900) xor estimated(901) xor estimated(902) xor estimated(903) xor estimated(904) xor estimated(905) xor estimated(906) xor estimated(907) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(912) xor estimated(913) xor estimated(914) xor estimated(915) xor estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(928) xor estimated(929) xor estimated(930) xor estimated(931) xor estimated(932) xor estimated(933) xor estimated(934) xor estimated(935) xor estimated(936) xor estimated(937) xor estimated(938) xor estimated(939) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(944) xor estimated(945) xor estimated(946) xor estimated(947) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(8) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(9) <= estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(10) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(11) <= estimated(800) xor estimated(801) xor estimated(802) xor estimated(803) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(12) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(13) <= estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(14) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(15) <= estimated(928) xor estimated(929) xor estimated(930) xor estimated(931) xor estimated(932) xor estimated(933) xor estimated(934) xor estimated(935) xor estimated(936) xor estimated(937) xor estimated(938) xor estimated(939) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(944) xor estimated(945) xor estimated(946) xor estimated(947) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(16) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(17) <= estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(18) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(19) <= estimated(784) xor estimated(785) xor estimated(786) xor estimated(787) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(20) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(21) <= estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(22) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(23) <= estimated(912) xor estimated(913) xor estimated(914) xor estimated(915) xor estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(944) xor estimated(945) xor estimated(946) xor estimated(947) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(24) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(25) <= estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(26) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(27) <= estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(28) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(29) <= estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(30) <= estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(31) <= estimated(944) xor estimated(945) xor estimated(946) xor estimated(947) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(32) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(33) <= estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(34) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(35) <= estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(36) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(37) <= estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(38) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(39) <= estimated(904) xor estimated(905) xor estimated(906) xor estimated(907) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(936) xor estimated(937) xor estimated(938) xor estimated(939) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(40) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(41) <= estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(42) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(43) <= estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(44) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(45) <= estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(46) <= estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(47) <= estimated(936) xor estimated(937) xor estimated(938) xor estimated(939) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(48) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(49) <= estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(50) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(51) <= estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(52) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(53) <= estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(54) <= estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(55) <= estimated(920) xor estimated(921) xor estimated(922) xor estimated(923) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(56) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(57) <= estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(58) <= estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(59) <= estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(60) <= estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(61) <= estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(62) <= estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(63) <= estimated(952) xor estimated(953) xor estimated(954) xor estimated(955) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(64) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(65) <= estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(66) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(67) <= estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(68) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(69) <= estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(70) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(71) <= estimated(900) xor estimated(901) xor estimated(902) xor estimated(903) xor estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(932) xor estimated(933) xor estimated(934) xor estimated(935) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(72) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(73) <= estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(74) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(75) <= estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(76) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(77) <= estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(78) <= estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(79) <= estimated(932) xor estimated(933) xor estimated(934) xor estimated(935) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(80) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(81) <= estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(82) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(83) <= estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(84) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(85) <= estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(86) <= estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(87) <= estimated(916) xor estimated(917) xor estimated(918) xor estimated(919) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(88) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(89) <= estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(90) <= estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(91) <= estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(92) <= estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(93) <= estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(94) <= estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(95) <= estimated(948) xor estimated(949) xor estimated(950) xor estimated(951) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(96) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(97) <= estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(98) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(99) <= estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(100) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(101) <= estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(102) <= estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(103) <= estimated(908) xor estimated(909) xor estimated(910) xor estimated(911) xor estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(104) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(105) <= estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(106) <= estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(107) <= estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(108) <= estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(109) <= estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(110) <= estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(111) <= estimated(940) xor estimated(941) xor estimated(942) xor estimated(943) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(112) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(113) <= estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(114) <= estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(115) <= estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(116) <= estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(117) <= estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(118) <= estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(119) <= estimated(924) xor estimated(925) xor estimated(926) xor estimated(927) xor estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(120) <= estimated(60) xor estimated(61) xor estimated(62) xor estimated(63);
partial_sums(7)(121) <= estimated(572) xor estimated(573) xor estimated(574) xor estimated(575);
partial_sums(7)(122) <= estimated(316) xor estimated(317) xor estimated(318) xor estimated(319);
partial_sums(7)(123) <= estimated(828) xor estimated(829) xor estimated(830) xor estimated(831);
partial_sums(7)(124) <= estimated(188) xor estimated(189) xor estimated(190) xor estimated(191);
partial_sums(7)(125) <= estimated(700) xor estimated(701) xor estimated(702) xor estimated(703);
partial_sums(7)(126) <= estimated(444) xor estimated(445) xor estimated(446) xor estimated(447);
partial_sums(7)(127) <= estimated(956) xor estimated(957) xor estimated(958) xor estimated(959);
partial_sums(7)(128) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(129) <= estimated(514) xor estimated(515) xor estimated(518) xor estimated(519) xor estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(546) xor estimated(547) xor estimated(550) xor estimated(551) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(130) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(131) <= estimated(770) xor estimated(771) xor estimated(774) xor estimated(775) xor estimated(778) xor estimated(779) xor estimated(782) xor estimated(783) xor estimated(786) xor estimated(787) xor estimated(790) xor estimated(791) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(802) xor estimated(803) xor estimated(806) xor estimated(807) xor estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(132) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(133) <= estimated(642) xor estimated(643) xor estimated(646) xor estimated(647) xor estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(674) xor estimated(675) xor estimated(678) xor estimated(679) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(134) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(135) <= estimated(898) xor estimated(899) xor estimated(902) xor estimated(903) xor estimated(906) xor estimated(907) xor estimated(910) xor estimated(911) xor estimated(914) xor estimated(915) xor estimated(918) xor estimated(919) xor estimated(922) xor estimated(923) xor estimated(926) xor estimated(927) xor estimated(930) xor estimated(931) xor estimated(934) xor estimated(935) xor estimated(938) xor estimated(939) xor estimated(942) xor estimated(943) xor estimated(946) xor estimated(947) xor estimated(950) xor estimated(951) xor estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(136) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(137) <= estimated(546) xor estimated(547) xor estimated(550) xor estimated(551) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(138) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(139) <= estimated(802) xor estimated(803) xor estimated(806) xor estimated(807) xor estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(140) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(141) <= estimated(674) xor estimated(675) xor estimated(678) xor estimated(679) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(142) <= estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(143) <= estimated(930) xor estimated(931) xor estimated(934) xor estimated(935) xor estimated(938) xor estimated(939) xor estimated(942) xor estimated(943) xor estimated(946) xor estimated(947) xor estimated(950) xor estimated(951) xor estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(144) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(145) <= estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(146) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(147) <= estimated(786) xor estimated(787) xor estimated(790) xor estimated(791) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(148) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(149) <= estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(150) <= estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(151) <= estimated(914) xor estimated(915) xor estimated(918) xor estimated(919) xor estimated(922) xor estimated(923) xor estimated(926) xor estimated(927) xor estimated(946) xor estimated(947) xor estimated(950) xor estimated(951) xor estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(152) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(153) <= estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(154) <= estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(155) <= estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(156) <= estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(157) <= estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(158) <= estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(159) <= estimated(946) xor estimated(947) xor estimated(950) xor estimated(951) xor estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(160) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(161) <= estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(162) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(163) <= estimated(778) xor estimated(779) xor estimated(782) xor estimated(783) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(164) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(165) <= estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(166) <= estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(167) <= estimated(906) xor estimated(907) xor estimated(910) xor estimated(911) xor estimated(922) xor estimated(923) xor estimated(926) xor estimated(927) xor estimated(938) xor estimated(939) xor estimated(942) xor estimated(943) xor estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(168) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(169) <= estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(170) <= estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(171) <= estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(172) <= estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(173) <= estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(174) <= estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(175) <= estimated(938) xor estimated(939) xor estimated(942) xor estimated(943) xor estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(176) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(177) <= estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(178) <= estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(179) <= estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(180) <= estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(181) <= estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(182) <= estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(183) <= estimated(922) xor estimated(923) xor estimated(926) xor estimated(927) xor estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(184) <= estimated(58) xor estimated(59) xor estimated(62) xor estimated(63);
partial_sums(7)(185) <= estimated(570) xor estimated(571) xor estimated(574) xor estimated(575);
partial_sums(7)(186) <= estimated(314) xor estimated(315) xor estimated(318) xor estimated(319);
partial_sums(7)(187) <= estimated(826) xor estimated(827) xor estimated(830) xor estimated(831);
partial_sums(7)(188) <= estimated(186) xor estimated(187) xor estimated(190) xor estimated(191);
partial_sums(7)(189) <= estimated(698) xor estimated(699) xor estimated(702) xor estimated(703);
partial_sums(7)(190) <= estimated(442) xor estimated(443) xor estimated(446) xor estimated(447);
partial_sums(7)(191) <= estimated(954) xor estimated(955) xor estimated(958) xor estimated(959);
partial_sums(7)(192) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(193) <= estimated(518) xor estimated(519) xor estimated(526) xor estimated(527) xor estimated(534) xor estimated(535) xor estimated(542) xor estimated(543) xor estimated(550) xor estimated(551) xor estimated(558) xor estimated(559) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575);
partial_sums(7)(194) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(195) <= estimated(774) xor estimated(775) xor estimated(782) xor estimated(783) xor estimated(790) xor estimated(791) xor estimated(798) xor estimated(799) xor estimated(806) xor estimated(807) xor estimated(814) xor estimated(815) xor estimated(822) xor estimated(823) xor estimated(830) xor estimated(831);
partial_sums(7)(196) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(197) <= estimated(646) xor estimated(647) xor estimated(654) xor estimated(655) xor estimated(662) xor estimated(663) xor estimated(670) xor estimated(671) xor estimated(678) xor estimated(679) xor estimated(686) xor estimated(687) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703);
partial_sums(7)(198) <= estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(199) <= estimated(902) xor estimated(903) xor estimated(910) xor estimated(911) xor estimated(918) xor estimated(919) xor estimated(926) xor estimated(927) xor estimated(934) xor estimated(935) xor estimated(942) xor estimated(943) xor estimated(950) xor estimated(951) xor estimated(958) xor estimated(959);
partial_sums(7)(200) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(201) <= estimated(550) xor estimated(551) xor estimated(558) xor estimated(559) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575);
partial_sums(7)(202) <= estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(203) <= estimated(806) xor estimated(807) xor estimated(814) xor estimated(815) xor estimated(822) xor estimated(823) xor estimated(830) xor estimated(831);
partial_sums(7)(204) <= estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(205) <= estimated(678) xor estimated(679) xor estimated(686) xor estimated(687) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703);
partial_sums(7)(206) <= estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(207) <= estimated(934) xor estimated(935) xor estimated(942) xor estimated(943) xor estimated(950) xor estimated(951) xor estimated(958) xor estimated(959);
partial_sums(7)(208) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(209) <= estimated(534) xor estimated(535) xor estimated(542) xor estimated(543) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575);
partial_sums(7)(210) <= estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(211) <= estimated(790) xor estimated(791) xor estimated(798) xor estimated(799) xor estimated(822) xor estimated(823) xor estimated(830) xor estimated(831);
partial_sums(7)(212) <= estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(213) <= estimated(662) xor estimated(663) xor estimated(670) xor estimated(671) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703);
partial_sums(7)(214) <= estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(215) <= estimated(918) xor estimated(919) xor estimated(926) xor estimated(927) xor estimated(950) xor estimated(951) xor estimated(958) xor estimated(959);
partial_sums(7)(216) <= estimated(54) xor estimated(55) xor estimated(62) xor estimated(63);
partial_sums(7)(217) <= estimated(566) xor estimated(567) xor estimated(574) xor estimated(575);
partial_sums(7)(218) <= estimated(310) xor estimated(311) xor estimated(318) xor estimated(319);
partial_sums(7)(219) <= estimated(822) xor estimated(823) xor estimated(830) xor estimated(831);
partial_sums(7)(220) <= estimated(182) xor estimated(183) xor estimated(190) xor estimated(191);
partial_sums(7)(221) <= estimated(694) xor estimated(695) xor estimated(702) xor estimated(703);
partial_sums(7)(222) <= estimated(438) xor estimated(439) xor estimated(446) xor estimated(447);
partial_sums(7)(223) <= estimated(950) xor estimated(951) xor estimated(958) xor estimated(959);
partial_sums(7)(224) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31) xor estimated(46) xor estimated(47) xor estimated(62) xor estimated(63);
partial_sums(7)(225) <= estimated(526) xor estimated(527) xor estimated(542) xor estimated(543) xor estimated(558) xor estimated(559) xor estimated(574) xor estimated(575);
partial_sums(7)(226) <= estimated(270) xor estimated(271) xor estimated(286) xor estimated(287) xor estimated(302) xor estimated(303) xor estimated(318) xor estimated(319);
partial_sums(7)(227) <= estimated(782) xor estimated(783) xor estimated(798) xor estimated(799) xor estimated(814) xor estimated(815) xor estimated(830) xor estimated(831);
partial_sums(7)(228) <= estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191);
partial_sums(7)(229) <= estimated(654) xor estimated(655) xor estimated(670) xor estimated(671) xor estimated(686) xor estimated(687) xor estimated(702) xor estimated(703);
partial_sums(7)(230) <= estimated(398) xor estimated(399) xor estimated(414) xor estimated(415) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447);
partial_sums(7)(231) <= estimated(910) xor estimated(911) xor estimated(926) xor estimated(927) xor estimated(942) xor estimated(943) xor estimated(958) xor estimated(959);
partial_sums(7)(232) <= estimated(46) xor estimated(47) xor estimated(62) xor estimated(63);
partial_sums(7)(233) <= estimated(558) xor estimated(559) xor estimated(574) xor estimated(575);
partial_sums(7)(234) <= estimated(302) xor estimated(303) xor estimated(318) xor estimated(319);
partial_sums(7)(235) <= estimated(814) xor estimated(815) xor estimated(830) xor estimated(831);
partial_sums(7)(236) <= estimated(174) xor estimated(175) xor estimated(190) xor estimated(191);
partial_sums(7)(237) <= estimated(686) xor estimated(687) xor estimated(702) xor estimated(703);
partial_sums(7)(238) <= estimated(430) xor estimated(431) xor estimated(446) xor estimated(447);
partial_sums(7)(239) <= estimated(942) xor estimated(943) xor estimated(958) xor estimated(959);
partial_sums(7)(240) <= estimated(30) xor estimated(31) xor estimated(62) xor estimated(63);
partial_sums(7)(241) <= estimated(542) xor estimated(543) xor estimated(574) xor estimated(575);
partial_sums(7)(242) <= estimated(286) xor estimated(287) xor estimated(318) xor estimated(319);
partial_sums(7)(243) <= estimated(798) xor estimated(799) xor estimated(830) xor estimated(831);
partial_sums(7)(244) <= estimated(158) xor estimated(159) xor estimated(190) xor estimated(191);
partial_sums(7)(245) <= estimated(670) xor estimated(671) xor estimated(702) xor estimated(703);
partial_sums(7)(246) <= estimated(414) xor estimated(415) xor estimated(446) xor estimated(447);
partial_sums(7)(247) <= estimated(926) xor estimated(927) xor estimated(958) xor estimated(959);
partial_sums(7)(248) <= estimated(62) xor estimated(63);
partial_sums(7)(249) <= estimated(574) xor estimated(575);
partial_sums(7)(250) <= estimated(318) xor estimated(319);
partial_sums(7)(251) <= estimated(830) xor estimated(831);
partial_sums(7)(252) <= estimated(190) xor estimated(191);
partial_sums(7)(253) <= estimated(702) xor estimated(703);
partial_sums(7)(254) <= estimated(446) xor estimated(447);
partial_sums(7)(255) <= estimated(958) xor estimated(959);
partial_sums(7)(256) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(257) <= estimated(513) xor estimated(515) xor estimated(517) xor estimated(519) xor estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(545) xor estimated(547) xor estimated(549) xor estimated(551) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(258) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(259) <= estimated(769) xor estimated(771) xor estimated(773) xor estimated(775) xor estimated(777) xor estimated(779) xor estimated(781) xor estimated(783) xor estimated(785) xor estimated(787) xor estimated(789) xor estimated(791) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(801) xor estimated(803) xor estimated(805) xor estimated(807) xor estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(260) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(261) <= estimated(641) xor estimated(643) xor estimated(645) xor estimated(647) xor estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(673) xor estimated(675) xor estimated(677) xor estimated(679) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(262) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(263) <= estimated(897) xor estimated(899) xor estimated(901) xor estimated(903) xor estimated(905) xor estimated(907) xor estimated(909) xor estimated(911) xor estimated(913) xor estimated(915) xor estimated(917) xor estimated(919) xor estimated(921) xor estimated(923) xor estimated(925) xor estimated(927) xor estimated(929) xor estimated(931) xor estimated(933) xor estimated(935) xor estimated(937) xor estimated(939) xor estimated(941) xor estimated(943) xor estimated(945) xor estimated(947) xor estimated(949) xor estimated(951) xor estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(264) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(265) <= estimated(545) xor estimated(547) xor estimated(549) xor estimated(551) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(266) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(267) <= estimated(801) xor estimated(803) xor estimated(805) xor estimated(807) xor estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(268) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(269) <= estimated(673) xor estimated(675) xor estimated(677) xor estimated(679) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(270) <= estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(271) <= estimated(929) xor estimated(931) xor estimated(933) xor estimated(935) xor estimated(937) xor estimated(939) xor estimated(941) xor estimated(943) xor estimated(945) xor estimated(947) xor estimated(949) xor estimated(951) xor estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(272) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(273) <= estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(274) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(275) <= estimated(785) xor estimated(787) xor estimated(789) xor estimated(791) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(276) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(277) <= estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(278) <= estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(279) <= estimated(913) xor estimated(915) xor estimated(917) xor estimated(919) xor estimated(921) xor estimated(923) xor estimated(925) xor estimated(927) xor estimated(945) xor estimated(947) xor estimated(949) xor estimated(951) xor estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(280) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(281) <= estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(282) <= estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(283) <= estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(284) <= estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(285) <= estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(286) <= estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(287) <= estimated(945) xor estimated(947) xor estimated(949) xor estimated(951) xor estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(288) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(289) <= estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(290) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(291) <= estimated(777) xor estimated(779) xor estimated(781) xor estimated(783) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(292) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(293) <= estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(294) <= estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(295) <= estimated(905) xor estimated(907) xor estimated(909) xor estimated(911) xor estimated(921) xor estimated(923) xor estimated(925) xor estimated(927) xor estimated(937) xor estimated(939) xor estimated(941) xor estimated(943) xor estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(296) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(297) <= estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(298) <= estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(299) <= estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(300) <= estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(301) <= estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(302) <= estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(303) <= estimated(937) xor estimated(939) xor estimated(941) xor estimated(943) xor estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(304) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(305) <= estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(306) <= estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(307) <= estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(308) <= estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(309) <= estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(310) <= estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(311) <= estimated(921) xor estimated(923) xor estimated(925) xor estimated(927) xor estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(312) <= estimated(57) xor estimated(59) xor estimated(61) xor estimated(63);
partial_sums(7)(313) <= estimated(569) xor estimated(571) xor estimated(573) xor estimated(575);
partial_sums(7)(314) <= estimated(313) xor estimated(315) xor estimated(317) xor estimated(319);
partial_sums(7)(315) <= estimated(825) xor estimated(827) xor estimated(829) xor estimated(831);
partial_sums(7)(316) <= estimated(185) xor estimated(187) xor estimated(189) xor estimated(191);
partial_sums(7)(317) <= estimated(697) xor estimated(699) xor estimated(701) xor estimated(703);
partial_sums(7)(318) <= estimated(441) xor estimated(443) xor estimated(445) xor estimated(447);
partial_sums(7)(319) <= estimated(953) xor estimated(955) xor estimated(957) xor estimated(959);
partial_sums(7)(320) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(321) <= estimated(517) xor estimated(519) xor estimated(525) xor estimated(527) xor estimated(533) xor estimated(535) xor estimated(541) xor estimated(543) xor estimated(549) xor estimated(551) xor estimated(557) xor estimated(559) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575);
partial_sums(7)(322) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(323) <= estimated(773) xor estimated(775) xor estimated(781) xor estimated(783) xor estimated(789) xor estimated(791) xor estimated(797) xor estimated(799) xor estimated(805) xor estimated(807) xor estimated(813) xor estimated(815) xor estimated(821) xor estimated(823) xor estimated(829) xor estimated(831);
partial_sums(7)(324) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(325) <= estimated(645) xor estimated(647) xor estimated(653) xor estimated(655) xor estimated(661) xor estimated(663) xor estimated(669) xor estimated(671) xor estimated(677) xor estimated(679) xor estimated(685) xor estimated(687) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703);
partial_sums(7)(326) <= estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(327) <= estimated(901) xor estimated(903) xor estimated(909) xor estimated(911) xor estimated(917) xor estimated(919) xor estimated(925) xor estimated(927) xor estimated(933) xor estimated(935) xor estimated(941) xor estimated(943) xor estimated(949) xor estimated(951) xor estimated(957) xor estimated(959);
partial_sums(7)(328) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(329) <= estimated(549) xor estimated(551) xor estimated(557) xor estimated(559) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575);
partial_sums(7)(330) <= estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(331) <= estimated(805) xor estimated(807) xor estimated(813) xor estimated(815) xor estimated(821) xor estimated(823) xor estimated(829) xor estimated(831);
partial_sums(7)(332) <= estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(333) <= estimated(677) xor estimated(679) xor estimated(685) xor estimated(687) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703);
partial_sums(7)(334) <= estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(335) <= estimated(933) xor estimated(935) xor estimated(941) xor estimated(943) xor estimated(949) xor estimated(951) xor estimated(957) xor estimated(959);
partial_sums(7)(336) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(337) <= estimated(533) xor estimated(535) xor estimated(541) xor estimated(543) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575);
partial_sums(7)(338) <= estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(339) <= estimated(789) xor estimated(791) xor estimated(797) xor estimated(799) xor estimated(821) xor estimated(823) xor estimated(829) xor estimated(831);
partial_sums(7)(340) <= estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(341) <= estimated(661) xor estimated(663) xor estimated(669) xor estimated(671) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703);
partial_sums(7)(342) <= estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(343) <= estimated(917) xor estimated(919) xor estimated(925) xor estimated(927) xor estimated(949) xor estimated(951) xor estimated(957) xor estimated(959);
partial_sums(7)(344) <= estimated(53) xor estimated(55) xor estimated(61) xor estimated(63);
partial_sums(7)(345) <= estimated(565) xor estimated(567) xor estimated(573) xor estimated(575);
partial_sums(7)(346) <= estimated(309) xor estimated(311) xor estimated(317) xor estimated(319);
partial_sums(7)(347) <= estimated(821) xor estimated(823) xor estimated(829) xor estimated(831);
partial_sums(7)(348) <= estimated(181) xor estimated(183) xor estimated(189) xor estimated(191);
partial_sums(7)(349) <= estimated(693) xor estimated(695) xor estimated(701) xor estimated(703);
partial_sums(7)(350) <= estimated(437) xor estimated(439) xor estimated(445) xor estimated(447);
partial_sums(7)(351) <= estimated(949) xor estimated(951) xor estimated(957) xor estimated(959);
partial_sums(7)(352) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31) xor estimated(45) xor estimated(47) xor estimated(61) xor estimated(63);
partial_sums(7)(353) <= estimated(525) xor estimated(527) xor estimated(541) xor estimated(543) xor estimated(557) xor estimated(559) xor estimated(573) xor estimated(575);
partial_sums(7)(354) <= estimated(269) xor estimated(271) xor estimated(285) xor estimated(287) xor estimated(301) xor estimated(303) xor estimated(317) xor estimated(319);
partial_sums(7)(355) <= estimated(781) xor estimated(783) xor estimated(797) xor estimated(799) xor estimated(813) xor estimated(815) xor estimated(829) xor estimated(831);
partial_sums(7)(356) <= estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191);
partial_sums(7)(357) <= estimated(653) xor estimated(655) xor estimated(669) xor estimated(671) xor estimated(685) xor estimated(687) xor estimated(701) xor estimated(703);
partial_sums(7)(358) <= estimated(397) xor estimated(399) xor estimated(413) xor estimated(415) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447);
partial_sums(7)(359) <= estimated(909) xor estimated(911) xor estimated(925) xor estimated(927) xor estimated(941) xor estimated(943) xor estimated(957) xor estimated(959);
partial_sums(7)(360) <= estimated(45) xor estimated(47) xor estimated(61) xor estimated(63);
partial_sums(7)(361) <= estimated(557) xor estimated(559) xor estimated(573) xor estimated(575);
partial_sums(7)(362) <= estimated(301) xor estimated(303) xor estimated(317) xor estimated(319);
partial_sums(7)(363) <= estimated(813) xor estimated(815) xor estimated(829) xor estimated(831);
partial_sums(7)(364) <= estimated(173) xor estimated(175) xor estimated(189) xor estimated(191);
partial_sums(7)(365) <= estimated(685) xor estimated(687) xor estimated(701) xor estimated(703);
partial_sums(7)(366) <= estimated(429) xor estimated(431) xor estimated(445) xor estimated(447);
partial_sums(7)(367) <= estimated(941) xor estimated(943) xor estimated(957) xor estimated(959);
partial_sums(7)(368) <= estimated(29) xor estimated(31) xor estimated(61) xor estimated(63);
partial_sums(7)(369) <= estimated(541) xor estimated(543) xor estimated(573) xor estimated(575);
partial_sums(7)(370) <= estimated(285) xor estimated(287) xor estimated(317) xor estimated(319);
partial_sums(7)(371) <= estimated(797) xor estimated(799) xor estimated(829) xor estimated(831);
partial_sums(7)(372) <= estimated(157) xor estimated(159) xor estimated(189) xor estimated(191);
partial_sums(7)(373) <= estimated(669) xor estimated(671) xor estimated(701) xor estimated(703);
partial_sums(7)(374) <= estimated(413) xor estimated(415) xor estimated(445) xor estimated(447);
partial_sums(7)(375) <= estimated(925) xor estimated(927) xor estimated(957) xor estimated(959);
partial_sums(7)(376) <= estimated(61) xor estimated(63);
partial_sums(7)(377) <= estimated(573) xor estimated(575);
partial_sums(7)(378) <= estimated(317) xor estimated(319);
partial_sums(7)(379) <= estimated(829) xor estimated(831);
partial_sums(7)(380) <= estimated(189) xor estimated(191);
partial_sums(7)(381) <= estimated(701) xor estimated(703);
partial_sums(7)(382) <= estimated(445) xor estimated(447);
partial_sums(7)(383) <= estimated(957) xor estimated(959);
partial_sums(7)(384) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(385) <= estimated(515) xor estimated(519) xor estimated(523) xor estimated(527) xor estimated(531) xor estimated(535) xor estimated(539) xor estimated(543) xor estimated(547) xor estimated(551) xor estimated(555) xor estimated(559) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575);
partial_sums(7)(386) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(387) <= estimated(771) xor estimated(775) xor estimated(779) xor estimated(783) xor estimated(787) xor estimated(791) xor estimated(795) xor estimated(799) xor estimated(803) xor estimated(807) xor estimated(811) xor estimated(815) xor estimated(819) xor estimated(823) xor estimated(827) xor estimated(831);
partial_sums(7)(388) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(389) <= estimated(643) xor estimated(647) xor estimated(651) xor estimated(655) xor estimated(659) xor estimated(663) xor estimated(667) xor estimated(671) xor estimated(675) xor estimated(679) xor estimated(683) xor estimated(687) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703);
partial_sums(7)(390) <= estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(391) <= estimated(899) xor estimated(903) xor estimated(907) xor estimated(911) xor estimated(915) xor estimated(919) xor estimated(923) xor estimated(927) xor estimated(931) xor estimated(935) xor estimated(939) xor estimated(943) xor estimated(947) xor estimated(951) xor estimated(955) xor estimated(959);
partial_sums(7)(392) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(393) <= estimated(547) xor estimated(551) xor estimated(555) xor estimated(559) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575);
partial_sums(7)(394) <= estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(395) <= estimated(803) xor estimated(807) xor estimated(811) xor estimated(815) xor estimated(819) xor estimated(823) xor estimated(827) xor estimated(831);
partial_sums(7)(396) <= estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(397) <= estimated(675) xor estimated(679) xor estimated(683) xor estimated(687) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703);
partial_sums(7)(398) <= estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(399) <= estimated(931) xor estimated(935) xor estimated(939) xor estimated(943) xor estimated(947) xor estimated(951) xor estimated(955) xor estimated(959);
partial_sums(7)(400) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(401) <= estimated(531) xor estimated(535) xor estimated(539) xor estimated(543) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575);
partial_sums(7)(402) <= estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(403) <= estimated(787) xor estimated(791) xor estimated(795) xor estimated(799) xor estimated(819) xor estimated(823) xor estimated(827) xor estimated(831);
partial_sums(7)(404) <= estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(405) <= estimated(659) xor estimated(663) xor estimated(667) xor estimated(671) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703);
partial_sums(7)(406) <= estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(407) <= estimated(915) xor estimated(919) xor estimated(923) xor estimated(927) xor estimated(947) xor estimated(951) xor estimated(955) xor estimated(959);
partial_sums(7)(408) <= estimated(51) xor estimated(55) xor estimated(59) xor estimated(63);
partial_sums(7)(409) <= estimated(563) xor estimated(567) xor estimated(571) xor estimated(575);
partial_sums(7)(410) <= estimated(307) xor estimated(311) xor estimated(315) xor estimated(319);
partial_sums(7)(411) <= estimated(819) xor estimated(823) xor estimated(827) xor estimated(831);
partial_sums(7)(412) <= estimated(179) xor estimated(183) xor estimated(187) xor estimated(191);
partial_sums(7)(413) <= estimated(691) xor estimated(695) xor estimated(699) xor estimated(703);
partial_sums(7)(414) <= estimated(435) xor estimated(439) xor estimated(443) xor estimated(447);
partial_sums(7)(415) <= estimated(947) xor estimated(951) xor estimated(955) xor estimated(959);
partial_sums(7)(416) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31) xor estimated(43) xor estimated(47) xor estimated(59) xor estimated(63);
partial_sums(7)(417) <= estimated(523) xor estimated(527) xor estimated(539) xor estimated(543) xor estimated(555) xor estimated(559) xor estimated(571) xor estimated(575);
partial_sums(7)(418) <= estimated(267) xor estimated(271) xor estimated(283) xor estimated(287) xor estimated(299) xor estimated(303) xor estimated(315) xor estimated(319);
partial_sums(7)(419) <= estimated(779) xor estimated(783) xor estimated(795) xor estimated(799) xor estimated(811) xor estimated(815) xor estimated(827) xor estimated(831);
partial_sums(7)(420) <= estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191);
partial_sums(7)(421) <= estimated(651) xor estimated(655) xor estimated(667) xor estimated(671) xor estimated(683) xor estimated(687) xor estimated(699) xor estimated(703);
partial_sums(7)(422) <= estimated(395) xor estimated(399) xor estimated(411) xor estimated(415) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447);
partial_sums(7)(423) <= estimated(907) xor estimated(911) xor estimated(923) xor estimated(927) xor estimated(939) xor estimated(943) xor estimated(955) xor estimated(959);
partial_sums(7)(424) <= estimated(43) xor estimated(47) xor estimated(59) xor estimated(63);
partial_sums(7)(425) <= estimated(555) xor estimated(559) xor estimated(571) xor estimated(575);
partial_sums(7)(426) <= estimated(299) xor estimated(303) xor estimated(315) xor estimated(319);
partial_sums(7)(427) <= estimated(811) xor estimated(815) xor estimated(827) xor estimated(831);
partial_sums(7)(428) <= estimated(171) xor estimated(175) xor estimated(187) xor estimated(191);
partial_sums(7)(429) <= estimated(683) xor estimated(687) xor estimated(699) xor estimated(703);
partial_sums(7)(430) <= estimated(427) xor estimated(431) xor estimated(443) xor estimated(447);
partial_sums(7)(431) <= estimated(939) xor estimated(943) xor estimated(955) xor estimated(959);
partial_sums(7)(432) <= estimated(27) xor estimated(31) xor estimated(59) xor estimated(63);
partial_sums(7)(433) <= estimated(539) xor estimated(543) xor estimated(571) xor estimated(575);
partial_sums(7)(434) <= estimated(283) xor estimated(287) xor estimated(315) xor estimated(319);
partial_sums(7)(435) <= estimated(795) xor estimated(799) xor estimated(827) xor estimated(831);
partial_sums(7)(436) <= estimated(155) xor estimated(159) xor estimated(187) xor estimated(191);
partial_sums(7)(437) <= estimated(667) xor estimated(671) xor estimated(699) xor estimated(703);
partial_sums(7)(438) <= estimated(411) xor estimated(415) xor estimated(443) xor estimated(447);
partial_sums(7)(439) <= estimated(923) xor estimated(927) xor estimated(955) xor estimated(959);
partial_sums(7)(440) <= estimated(59) xor estimated(63);
partial_sums(7)(441) <= estimated(571) xor estimated(575);
partial_sums(7)(442) <= estimated(315) xor estimated(319);
partial_sums(7)(443) <= estimated(827) xor estimated(831);
partial_sums(7)(444) <= estimated(187) xor estimated(191);
partial_sums(7)(445) <= estimated(699) xor estimated(703);
partial_sums(7)(446) <= estimated(443) xor estimated(447);
partial_sums(7)(447) <= estimated(955) xor estimated(959);
partial_sums(7)(448) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31) xor estimated(39) xor estimated(47) xor estimated(55) xor estimated(63);
partial_sums(7)(449) <= estimated(519) xor estimated(527) xor estimated(535) xor estimated(543) xor estimated(551) xor estimated(559) xor estimated(567) xor estimated(575);
partial_sums(7)(450) <= estimated(263) xor estimated(271) xor estimated(279) xor estimated(287) xor estimated(295) xor estimated(303) xor estimated(311) xor estimated(319);
partial_sums(7)(451) <= estimated(775) xor estimated(783) xor estimated(791) xor estimated(799) xor estimated(807) xor estimated(815) xor estimated(823) xor estimated(831);
partial_sums(7)(452) <= estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191);
partial_sums(7)(453) <= estimated(647) xor estimated(655) xor estimated(663) xor estimated(671) xor estimated(679) xor estimated(687) xor estimated(695) xor estimated(703);
partial_sums(7)(454) <= estimated(391) xor estimated(399) xor estimated(407) xor estimated(415) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447);
partial_sums(7)(455) <= estimated(903) xor estimated(911) xor estimated(919) xor estimated(927) xor estimated(935) xor estimated(943) xor estimated(951) xor estimated(959);
partial_sums(7)(456) <= estimated(39) xor estimated(47) xor estimated(55) xor estimated(63);
partial_sums(7)(457) <= estimated(551) xor estimated(559) xor estimated(567) xor estimated(575);
partial_sums(7)(458) <= estimated(295) xor estimated(303) xor estimated(311) xor estimated(319);
partial_sums(7)(459) <= estimated(807) xor estimated(815) xor estimated(823) xor estimated(831);
partial_sums(7)(460) <= estimated(167) xor estimated(175) xor estimated(183) xor estimated(191);
partial_sums(7)(461) <= estimated(679) xor estimated(687) xor estimated(695) xor estimated(703);
partial_sums(7)(462) <= estimated(423) xor estimated(431) xor estimated(439) xor estimated(447);
partial_sums(7)(463) <= estimated(935) xor estimated(943) xor estimated(951) xor estimated(959);
partial_sums(7)(464) <= estimated(23) xor estimated(31) xor estimated(55) xor estimated(63);
partial_sums(7)(465) <= estimated(535) xor estimated(543) xor estimated(567) xor estimated(575);
partial_sums(7)(466) <= estimated(279) xor estimated(287) xor estimated(311) xor estimated(319);
partial_sums(7)(467) <= estimated(791) xor estimated(799) xor estimated(823) xor estimated(831);
partial_sums(7)(468) <= estimated(151) xor estimated(159) xor estimated(183) xor estimated(191);
partial_sums(7)(469) <= estimated(663) xor estimated(671) xor estimated(695) xor estimated(703);
partial_sums(7)(470) <= estimated(407) xor estimated(415) xor estimated(439) xor estimated(447);
partial_sums(7)(471) <= estimated(919) xor estimated(927) xor estimated(951) xor estimated(959);
partial_sums(7)(472) <= estimated(55) xor estimated(63);
partial_sums(7)(473) <= estimated(567) xor estimated(575);
partial_sums(7)(474) <= estimated(311) xor estimated(319);
partial_sums(7)(475) <= estimated(823) xor estimated(831);
partial_sums(7)(476) <= estimated(183) xor estimated(191);
partial_sums(7)(477) <= estimated(695) xor estimated(703);
partial_sums(7)(478) <= estimated(439) xor estimated(447);
partial_sums(7)(479) <= estimated(951) xor estimated(959);
partial_sums(7)(480) <= estimated(15) xor estimated(31) xor estimated(47) xor estimated(63);
partial_sums(7)(481) <= estimated(527) xor estimated(543) xor estimated(559) xor estimated(575);
partial_sums(7)(482) <= estimated(271) xor estimated(287) xor estimated(303) xor estimated(319);
partial_sums(7)(483) <= estimated(783) xor estimated(799) xor estimated(815) xor estimated(831);
partial_sums(7)(484) <= estimated(143) xor estimated(159) xor estimated(175) xor estimated(191);
partial_sums(7)(485) <= estimated(655) xor estimated(671) xor estimated(687) xor estimated(703);
partial_sums(7)(486) <= estimated(399) xor estimated(415) xor estimated(431) xor estimated(447);
partial_sums(7)(487) <= estimated(911) xor estimated(927) xor estimated(943) xor estimated(959);
partial_sums(7)(488) <= estimated(47) xor estimated(63);
partial_sums(7)(489) <= estimated(559) xor estimated(575);
partial_sums(7)(490) <= estimated(303) xor estimated(319);
partial_sums(7)(491) <= estimated(815) xor estimated(831);
partial_sums(7)(492) <= estimated(175) xor estimated(191);
partial_sums(7)(493) <= estimated(687) xor estimated(703);
partial_sums(7)(494) <= estimated(431) xor estimated(447);
partial_sums(7)(495) <= estimated(943) xor estimated(959);
partial_sums(7)(496) <= estimated(31) xor estimated(63);
partial_sums(7)(497) <= estimated(543) xor estimated(575);
partial_sums(7)(498) <= estimated(287) xor estimated(319);
partial_sums(7)(499) <= estimated(799) xor estimated(831);
partial_sums(7)(500) <= estimated(159) xor estimated(191);
partial_sums(7)(501) <= estimated(671) xor estimated(703);
partial_sums(7)(502) <= estimated(415) xor estimated(447);
partial_sums(7)(503) <= estimated(927) xor estimated(959);
partial_sums(7)(504) <= estimated(63);
partial_sums(7)(505) <= estimated(575);
partial_sums(7)(506) <= estimated(319);
partial_sums(7)(507) <= estimated(831);
partial_sums(7)(508) <= estimated(191);
partial_sums(7)(509) <= estimated(703);
partial_sums(7)(510) <= estimated(447);
partial_sums(7)(511) <= estimated(959);
partial_sums(8)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(1) <= estimated(512) xor estimated(513) xor estimated(514) xor estimated(515) xor estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(576) xor estimated(577) xor estimated(578) xor estimated(579) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(2) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(3) <= estimated(768) xor estimated(769) xor estimated(770) xor estimated(771) xor estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(784) xor estimated(785) xor estimated(786) xor estimated(787) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(800) xor estimated(801) xor estimated(802) xor estimated(803) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(832) xor estimated(833) xor estimated(834) xor estimated(835) xor estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(848) xor estimated(849) xor estimated(850) xor estimated(851) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(864) xor estimated(865) xor estimated(866) xor estimated(867) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(4) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(5) <= estimated(576) xor estimated(577) xor estimated(578) xor estimated(579) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(6) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(7) <= estimated(832) xor estimated(833) xor estimated(834) xor estimated(835) xor estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(848) xor estimated(849) xor estimated(850) xor estimated(851) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(864) xor estimated(865) xor estimated(866) xor estimated(867) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(8) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(9) <= estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(10) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(11) <= estimated(800) xor estimated(801) xor estimated(802) xor estimated(803) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(864) xor estimated(865) xor estimated(866) xor estimated(867) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(12) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(13) <= estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(14) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(15) <= estimated(864) xor estimated(865) xor estimated(866) xor estimated(867) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(16) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(17) <= estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(18) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(19) <= estimated(784) xor estimated(785) xor estimated(786) xor estimated(787) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(848) xor estimated(849) xor estimated(850) xor estimated(851) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(20) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(21) <= estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(22) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(23) <= estimated(848) xor estimated(849) xor estimated(850) xor estimated(851) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(24) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(25) <= estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(26) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(27) <= estimated(816) xor estimated(817) xor estimated(818) xor estimated(819) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(28) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(29) <= estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(30) <= estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(31) <= estimated(880) xor estimated(881) xor estimated(882) xor estimated(883) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(32) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(33) <= estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(34) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(35) <= estimated(776) xor estimated(777) xor estimated(778) xor estimated(779) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(36) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(37) <= estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(38) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(39) <= estimated(840) xor estimated(841) xor estimated(842) xor estimated(843) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(40) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(41) <= estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(42) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(43) <= estimated(808) xor estimated(809) xor estimated(810) xor estimated(811) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(44) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(45) <= estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(46) <= estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(47) <= estimated(872) xor estimated(873) xor estimated(874) xor estimated(875) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(48) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(49) <= estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(50) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(51) <= estimated(792) xor estimated(793) xor estimated(794) xor estimated(795) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(52) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(53) <= estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(54) <= estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(55) <= estimated(856) xor estimated(857) xor estimated(858) xor estimated(859) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(56) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(57) <= estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(58) <= estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(59) <= estimated(824) xor estimated(825) xor estimated(826) xor estimated(827) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(60) <= estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(61) <= estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(62) <= estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(63) <= estimated(888) xor estimated(889) xor estimated(890) xor estimated(891) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(64) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(65) <= estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(66) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(67) <= estimated(772) xor estimated(773) xor estimated(774) xor estimated(775) xor estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(68) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(69) <= estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(70) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(71) <= estimated(836) xor estimated(837) xor estimated(838) xor estimated(839) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(72) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(73) <= estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(74) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(75) <= estimated(804) xor estimated(805) xor estimated(806) xor estimated(807) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(76) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(77) <= estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(78) <= estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(79) <= estimated(868) xor estimated(869) xor estimated(870) xor estimated(871) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(80) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(81) <= estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(82) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(83) <= estimated(788) xor estimated(789) xor estimated(790) xor estimated(791) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(84) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(85) <= estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(86) <= estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(87) <= estimated(852) xor estimated(853) xor estimated(854) xor estimated(855) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(88) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(89) <= estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(90) <= estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(91) <= estimated(820) xor estimated(821) xor estimated(822) xor estimated(823) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(92) <= estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(93) <= estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(94) <= estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(95) <= estimated(884) xor estimated(885) xor estimated(886) xor estimated(887) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(96) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(97) <= estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(98) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(99) <= estimated(780) xor estimated(781) xor estimated(782) xor estimated(783) xor estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(100) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(101) <= estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(102) <= estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(103) <= estimated(844) xor estimated(845) xor estimated(846) xor estimated(847) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(104) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(105) <= estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(106) <= estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(107) <= estimated(812) xor estimated(813) xor estimated(814) xor estimated(815) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(108) <= estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(109) <= estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(110) <= estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(111) <= estimated(876) xor estimated(877) xor estimated(878) xor estimated(879) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(112) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(113) <= estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(114) <= estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(115) <= estimated(796) xor estimated(797) xor estimated(798) xor estimated(799) xor estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(116) <= estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(117) <= estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(118) <= estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(119) <= estimated(860) xor estimated(861) xor estimated(862) xor estimated(863) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(120) <= estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(121) <= estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(122) <= estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(123) <= estimated(828) xor estimated(829) xor estimated(830) xor estimated(831) xor estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(124) <= estimated(124) xor estimated(125) xor estimated(126) xor estimated(127);
partial_sums(8)(125) <= estimated(636) xor estimated(637) xor estimated(638) xor estimated(639);
partial_sums(8)(126) <= estimated(380) xor estimated(381) xor estimated(382) xor estimated(383);
partial_sums(8)(127) <= estimated(892) xor estimated(893) xor estimated(894) xor estimated(895);
partial_sums(8)(128) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(129) <= estimated(514) xor estimated(515) xor estimated(518) xor estimated(519) xor estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(546) xor estimated(547) xor estimated(550) xor estimated(551) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(578) xor estimated(579) xor estimated(582) xor estimated(583) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(130) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(131) <= estimated(770) xor estimated(771) xor estimated(774) xor estimated(775) xor estimated(778) xor estimated(779) xor estimated(782) xor estimated(783) xor estimated(786) xor estimated(787) xor estimated(790) xor estimated(791) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(802) xor estimated(803) xor estimated(806) xor estimated(807) xor estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(834) xor estimated(835) xor estimated(838) xor estimated(839) xor estimated(842) xor estimated(843) xor estimated(846) xor estimated(847) xor estimated(850) xor estimated(851) xor estimated(854) xor estimated(855) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(866) xor estimated(867) xor estimated(870) xor estimated(871) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(132) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(133) <= estimated(578) xor estimated(579) xor estimated(582) xor estimated(583) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(134) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(135) <= estimated(834) xor estimated(835) xor estimated(838) xor estimated(839) xor estimated(842) xor estimated(843) xor estimated(846) xor estimated(847) xor estimated(850) xor estimated(851) xor estimated(854) xor estimated(855) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(866) xor estimated(867) xor estimated(870) xor estimated(871) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(136) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(137) <= estimated(546) xor estimated(547) xor estimated(550) xor estimated(551) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(138) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(139) <= estimated(802) xor estimated(803) xor estimated(806) xor estimated(807) xor estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(866) xor estimated(867) xor estimated(870) xor estimated(871) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(140) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(141) <= estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(142) <= estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(143) <= estimated(866) xor estimated(867) xor estimated(870) xor estimated(871) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(144) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(145) <= estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(146) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(147) <= estimated(786) xor estimated(787) xor estimated(790) xor estimated(791) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(850) xor estimated(851) xor estimated(854) xor estimated(855) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(148) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(149) <= estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(150) <= estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(151) <= estimated(850) xor estimated(851) xor estimated(854) xor estimated(855) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(152) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(153) <= estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(154) <= estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(155) <= estimated(818) xor estimated(819) xor estimated(822) xor estimated(823) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(156) <= estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(157) <= estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(158) <= estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(159) <= estimated(882) xor estimated(883) xor estimated(886) xor estimated(887) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(160) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(161) <= estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(162) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(163) <= estimated(778) xor estimated(779) xor estimated(782) xor estimated(783) xor estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(842) xor estimated(843) xor estimated(846) xor estimated(847) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(164) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(165) <= estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(166) <= estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(167) <= estimated(842) xor estimated(843) xor estimated(846) xor estimated(847) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(168) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(169) <= estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(170) <= estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(171) <= estimated(810) xor estimated(811) xor estimated(814) xor estimated(815) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(172) <= estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(173) <= estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(174) <= estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(175) <= estimated(874) xor estimated(875) xor estimated(878) xor estimated(879) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(176) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(177) <= estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(178) <= estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(179) <= estimated(794) xor estimated(795) xor estimated(798) xor estimated(799) xor estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(180) <= estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(181) <= estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(182) <= estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(183) <= estimated(858) xor estimated(859) xor estimated(862) xor estimated(863) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(184) <= estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(185) <= estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(186) <= estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(187) <= estimated(826) xor estimated(827) xor estimated(830) xor estimated(831) xor estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(188) <= estimated(122) xor estimated(123) xor estimated(126) xor estimated(127);
partial_sums(8)(189) <= estimated(634) xor estimated(635) xor estimated(638) xor estimated(639);
partial_sums(8)(190) <= estimated(378) xor estimated(379) xor estimated(382) xor estimated(383);
partial_sums(8)(191) <= estimated(890) xor estimated(891) xor estimated(894) xor estimated(895);
partial_sums(8)(192) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(193) <= estimated(518) xor estimated(519) xor estimated(526) xor estimated(527) xor estimated(534) xor estimated(535) xor estimated(542) xor estimated(543) xor estimated(550) xor estimated(551) xor estimated(558) xor estimated(559) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(582) xor estimated(583) xor estimated(590) xor estimated(591) xor estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(194) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(195) <= estimated(774) xor estimated(775) xor estimated(782) xor estimated(783) xor estimated(790) xor estimated(791) xor estimated(798) xor estimated(799) xor estimated(806) xor estimated(807) xor estimated(814) xor estimated(815) xor estimated(822) xor estimated(823) xor estimated(830) xor estimated(831) xor estimated(838) xor estimated(839) xor estimated(846) xor estimated(847) xor estimated(854) xor estimated(855) xor estimated(862) xor estimated(863) xor estimated(870) xor estimated(871) xor estimated(878) xor estimated(879) xor estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(196) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(197) <= estimated(582) xor estimated(583) xor estimated(590) xor estimated(591) xor estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(198) <= estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(199) <= estimated(838) xor estimated(839) xor estimated(846) xor estimated(847) xor estimated(854) xor estimated(855) xor estimated(862) xor estimated(863) xor estimated(870) xor estimated(871) xor estimated(878) xor estimated(879) xor estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(200) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(201) <= estimated(550) xor estimated(551) xor estimated(558) xor estimated(559) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(202) <= estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(203) <= estimated(806) xor estimated(807) xor estimated(814) xor estimated(815) xor estimated(822) xor estimated(823) xor estimated(830) xor estimated(831) xor estimated(870) xor estimated(871) xor estimated(878) xor estimated(879) xor estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(204) <= estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(205) <= estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(206) <= estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(207) <= estimated(870) xor estimated(871) xor estimated(878) xor estimated(879) xor estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(208) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(209) <= estimated(534) xor estimated(535) xor estimated(542) xor estimated(543) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(210) <= estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(211) <= estimated(790) xor estimated(791) xor estimated(798) xor estimated(799) xor estimated(822) xor estimated(823) xor estimated(830) xor estimated(831) xor estimated(854) xor estimated(855) xor estimated(862) xor estimated(863) xor estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(212) <= estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(213) <= estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(214) <= estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(215) <= estimated(854) xor estimated(855) xor estimated(862) xor estimated(863) xor estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(216) <= estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(217) <= estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(218) <= estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(219) <= estimated(822) xor estimated(823) xor estimated(830) xor estimated(831) xor estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(220) <= estimated(118) xor estimated(119) xor estimated(126) xor estimated(127);
partial_sums(8)(221) <= estimated(630) xor estimated(631) xor estimated(638) xor estimated(639);
partial_sums(8)(222) <= estimated(374) xor estimated(375) xor estimated(382) xor estimated(383);
partial_sums(8)(223) <= estimated(886) xor estimated(887) xor estimated(894) xor estimated(895);
partial_sums(8)(224) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31) xor estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(225) <= estimated(526) xor estimated(527) xor estimated(542) xor estimated(543) xor estimated(558) xor estimated(559) xor estimated(574) xor estimated(575) xor estimated(590) xor estimated(591) xor estimated(606) xor estimated(607) xor estimated(622) xor estimated(623) xor estimated(638) xor estimated(639);
partial_sums(8)(226) <= estimated(270) xor estimated(271) xor estimated(286) xor estimated(287) xor estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(227) <= estimated(782) xor estimated(783) xor estimated(798) xor estimated(799) xor estimated(814) xor estimated(815) xor estimated(830) xor estimated(831) xor estimated(846) xor estimated(847) xor estimated(862) xor estimated(863) xor estimated(878) xor estimated(879) xor estimated(894) xor estimated(895);
partial_sums(8)(228) <= estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(229) <= estimated(590) xor estimated(591) xor estimated(606) xor estimated(607) xor estimated(622) xor estimated(623) xor estimated(638) xor estimated(639);
partial_sums(8)(230) <= estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(231) <= estimated(846) xor estimated(847) xor estimated(862) xor estimated(863) xor estimated(878) xor estimated(879) xor estimated(894) xor estimated(895);
partial_sums(8)(232) <= estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(233) <= estimated(558) xor estimated(559) xor estimated(574) xor estimated(575) xor estimated(622) xor estimated(623) xor estimated(638) xor estimated(639);
partial_sums(8)(234) <= estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(235) <= estimated(814) xor estimated(815) xor estimated(830) xor estimated(831) xor estimated(878) xor estimated(879) xor estimated(894) xor estimated(895);
partial_sums(8)(236) <= estimated(110) xor estimated(111) xor estimated(126) xor estimated(127);
partial_sums(8)(237) <= estimated(622) xor estimated(623) xor estimated(638) xor estimated(639);
partial_sums(8)(238) <= estimated(366) xor estimated(367) xor estimated(382) xor estimated(383);
partial_sums(8)(239) <= estimated(878) xor estimated(879) xor estimated(894) xor estimated(895);
partial_sums(8)(240) <= estimated(30) xor estimated(31) xor estimated(62) xor estimated(63) xor estimated(94) xor estimated(95) xor estimated(126) xor estimated(127);
partial_sums(8)(241) <= estimated(542) xor estimated(543) xor estimated(574) xor estimated(575) xor estimated(606) xor estimated(607) xor estimated(638) xor estimated(639);
partial_sums(8)(242) <= estimated(286) xor estimated(287) xor estimated(318) xor estimated(319) xor estimated(350) xor estimated(351) xor estimated(382) xor estimated(383);
partial_sums(8)(243) <= estimated(798) xor estimated(799) xor estimated(830) xor estimated(831) xor estimated(862) xor estimated(863) xor estimated(894) xor estimated(895);
partial_sums(8)(244) <= estimated(94) xor estimated(95) xor estimated(126) xor estimated(127);
partial_sums(8)(245) <= estimated(606) xor estimated(607) xor estimated(638) xor estimated(639);
partial_sums(8)(246) <= estimated(350) xor estimated(351) xor estimated(382) xor estimated(383);
partial_sums(8)(247) <= estimated(862) xor estimated(863) xor estimated(894) xor estimated(895);
partial_sums(8)(248) <= estimated(62) xor estimated(63) xor estimated(126) xor estimated(127);
partial_sums(8)(249) <= estimated(574) xor estimated(575) xor estimated(638) xor estimated(639);
partial_sums(8)(250) <= estimated(318) xor estimated(319) xor estimated(382) xor estimated(383);
partial_sums(8)(251) <= estimated(830) xor estimated(831) xor estimated(894) xor estimated(895);
partial_sums(8)(252) <= estimated(126) xor estimated(127);
partial_sums(8)(253) <= estimated(638) xor estimated(639);
partial_sums(8)(254) <= estimated(382) xor estimated(383);
partial_sums(8)(255) <= estimated(894) xor estimated(895);
partial_sums(8)(256) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(257) <= estimated(513) xor estimated(515) xor estimated(517) xor estimated(519) xor estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(545) xor estimated(547) xor estimated(549) xor estimated(551) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(577) xor estimated(579) xor estimated(581) xor estimated(583) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(258) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(259) <= estimated(769) xor estimated(771) xor estimated(773) xor estimated(775) xor estimated(777) xor estimated(779) xor estimated(781) xor estimated(783) xor estimated(785) xor estimated(787) xor estimated(789) xor estimated(791) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(801) xor estimated(803) xor estimated(805) xor estimated(807) xor estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(833) xor estimated(835) xor estimated(837) xor estimated(839) xor estimated(841) xor estimated(843) xor estimated(845) xor estimated(847) xor estimated(849) xor estimated(851) xor estimated(853) xor estimated(855) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(865) xor estimated(867) xor estimated(869) xor estimated(871) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(260) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(261) <= estimated(577) xor estimated(579) xor estimated(581) xor estimated(583) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(262) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(263) <= estimated(833) xor estimated(835) xor estimated(837) xor estimated(839) xor estimated(841) xor estimated(843) xor estimated(845) xor estimated(847) xor estimated(849) xor estimated(851) xor estimated(853) xor estimated(855) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(865) xor estimated(867) xor estimated(869) xor estimated(871) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(264) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(265) <= estimated(545) xor estimated(547) xor estimated(549) xor estimated(551) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(266) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(267) <= estimated(801) xor estimated(803) xor estimated(805) xor estimated(807) xor estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(865) xor estimated(867) xor estimated(869) xor estimated(871) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(268) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(269) <= estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(270) <= estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(271) <= estimated(865) xor estimated(867) xor estimated(869) xor estimated(871) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(272) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(273) <= estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(274) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(275) <= estimated(785) xor estimated(787) xor estimated(789) xor estimated(791) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(849) xor estimated(851) xor estimated(853) xor estimated(855) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(276) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(277) <= estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(278) <= estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(279) <= estimated(849) xor estimated(851) xor estimated(853) xor estimated(855) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(280) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(281) <= estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(282) <= estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(283) <= estimated(817) xor estimated(819) xor estimated(821) xor estimated(823) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(284) <= estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(285) <= estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(286) <= estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(287) <= estimated(881) xor estimated(883) xor estimated(885) xor estimated(887) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(288) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(289) <= estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(290) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(291) <= estimated(777) xor estimated(779) xor estimated(781) xor estimated(783) xor estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(841) xor estimated(843) xor estimated(845) xor estimated(847) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(292) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(293) <= estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(294) <= estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(295) <= estimated(841) xor estimated(843) xor estimated(845) xor estimated(847) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(296) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(297) <= estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(298) <= estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(299) <= estimated(809) xor estimated(811) xor estimated(813) xor estimated(815) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(300) <= estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(301) <= estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(302) <= estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(303) <= estimated(873) xor estimated(875) xor estimated(877) xor estimated(879) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(304) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(305) <= estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(306) <= estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(307) <= estimated(793) xor estimated(795) xor estimated(797) xor estimated(799) xor estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(308) <= estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(309) <= estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(310) <= estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(311) <= estimated(857) xor estimated(859) xor estimated(861) xor estimated(863) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(312) <= estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(313) <= estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(314) <= estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(315) <= estimated(825) xor estimated(827) xor estimated(829) xor estimated(831) xor estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(316) <= estimated(121) xor estimated(123) xor estimated(125) xor estimated(127);
partial_sums(8)(317) <= estimated(633) xor estimated(635) xor estimated(637) xor estimated(639);
partial_sums(8)(318) <= estimated(377) xor estimated(379) xor estimated(381) xor estimated(383);
partial_sums(8)(319) <= estimated(889) xor estimated(891) xor estimated(893) xor estimated(895);
partial_sums(8)(320) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(321) <= estimated(517) xor estimated(519) xor estimated(525) xor estimated(527) xor estimated(533) xor estimated(535) xor estimated(541) xor estimated(543) xor estimated(549) xor estimated(551) xor estimated(557) xor estimated(559) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(581) xor estimated(583) xor estimated(589) xor estimated(591) xor estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(322) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(323) <= estimated(773) xor estimated(775) xor estimated(781) xor estimated(783) xor estimated(789) xor estimated(791) xor estimated(797) xor estimated(799) xor estimated(805) xor estimated(807) xor estimated(813) xor estimated(815) xor estimated(821) xor estimated(823) xor estimated(829) xor estimated(831) xor estimated(837) xor estimated(839) xor estimated(845) xor estimated(847) xor estimated(853) xor estimated(855) xor estimated(861) xor estimated(863) xor estimated(869) xor estimated(871) xor estimated(877) xor estimated(879) xor estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(324) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(325) <= estimated(581) xor estimated(583) xor estimated(589) xor estimated(591) xor estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(326) <= estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(327) <= estimated(837) xor estimated(839) xor estimated(845) xor estimated(847) xor estimated(853) xor estimated(855) xor estimated(861) xor estimated(863) xor estimated(869) xor estimated(871) xor estimated(877) xor estimated(879) xor estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(328) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(329) <= estimated(549) xor estimated(551) xor estimated(557) xor estimated(559) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(330) <= estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(331) <= estimated(805) xor estimated(807) xor estimated(813) xor estimated(815) xor estimated(821) xor estimated(823) xor estimated(829) xor estimated(831) xor estimated(869) xor estimated(871) xor estimated(877) xor estimated(879) xor estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(332) <= estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(333) <= estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(334) <= estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(335) <= estimated(869) xor estimated(871) xor estimated(877) xor estimated(879) xor estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(336) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(337) <= estimated(533) xor estimated(535) xor estimated(541) xor estimated(543) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(338) <= estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(339) <= estimated(789) xor estimated(791) xor estimated(797) xor estimated(799) xor estimated(821) xor estimated(823) xor estimated(829) xor estimated(831) xor estimated(853) xor estimated(855) xor estimated(861) xor estimated(863) xor estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(340) <= estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(341) <= estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(342) <= estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(343) <= estimated(853) xor estimated(855) xor estimated(861) xor estimated(863) xor estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(344) <= estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(345) <= estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(346) <= estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(347) <= estimated(821) xor estimated(823) xor estimated(829) xor estimated(831) xor estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(348) <= estimated(117) xor estimated(119) xor estimated(125) xor estimated(127);
partial_sums(8)(349) <= estimated(629) xor estimated(631) xor estimated(637) xor estimated(639);
partial_sums(8)(350) <= estimated(373) xor estimated(375) xor estimated(381) xor estimated(383);
partial_sums(8)(351) <= estimated(885) xor estimated(887) xor estimated(893) xor estimated(895);
partial_sums(8)(352) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31) xor estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(353) <= estimated(525) xor estimated(527) xor estimated(541) xor estimated(543) xor estimated(557) xor estimated(559) xor estimated(573) xor estimated(575) xor estimated(589) xor estimated(591) xor estimated(605) xor estimated(607) xor estimated(621) xor estimated(623) xor estimated(637) xor estimated(639);
partial_sums(8)(354) <= estimated(269) xor estimated(271) xor estimated(285) xor estimated(287) xor estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(355) <= estimated(781) xor estimated(783) xor estimated(797) xor estimated(799) xor estimated(813) xor estimated(815) xor estimated(829) xor estimated(831) xor estimated(845) xor estimated(847) xor estimated(861) xor estimated(863) xor estimated(877) xor estimated(879) xor estimated(893) xor estimated(895);
partial_sums(8)(356) <= estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(357) <= estimated(589) xor estimated(591) xor estimated(605) xor estimated(607) xor estimated(621) xor estimated(623) xor estimated(637) xor estimated(639);
partial_sums(8)(358) <= estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(359) <= estimated(845) xor estimated(847) xor estimated(861) xor estimated(863) xor estimated(877) xor estimated(879) xor estimated(893) xor estimated(895);
partial_sums(8)(360) <= estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(361) <= estimated(557) xor estimated(559) xor estimated(573) xor estimated(575) xor estimated(621) xor estimated(623) xor estimated(637) xor estimated(639);
partial_sums(8)(362) <= estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(363) <= estimated(813) xor estimated(815) xor estimated(829) xor estimated(831) xor estimated(877) xor estimated(879) xor estimated(893) xor estimated(895);
partial_sums(8)(364) <= estimated(109) xor estimated(111) xor estimated(125) xor estimated(127);
partial_sums(8)(365) <= estimated(621) xor estimated(623) xor estimated(637) xor estimated(639);
partial_sums(8)(366) <= estimated(365) xor estimated(367) xor estimated(381) xor estimated(383);
partial_sums(8)(367) <= estimated(877) xor estimated(879) xor estimated(893) xor estimated(895);
partial_sums(8)(368) <= estimated(29) xor estimated(31) xor estimated(61) xor estimated(63) xor estimated(93) xor estimated(95) xor estimated(125) xor estimated(127);
partial_sums(8)(369) <= estimated(541) xor estimated(543) xor estimated(573) xor estimated(575) xor estimated(605) xor estimated(607) xor estimated(637) xor estimated(639);
partial_sums(8)(370) <= estimated(285) xor estimated(287) xor estimated(317) xor estimated(319) xor estimated(349) xor estimated(351) xor estimated(381) xor estimated(383);
partial_sums(8)(371) <= estimated(797) xor estimated(799) xor estimated(829) xor estimated(831) xor estimated(861) xor estimated(863) xor estimated(893) xor estimated(895);
partial_sums(8)(372) <= estimated(93) xor estimated(95) xor estimated(125) xor estimated(127);
partial_sums(8)(373) <= estimated(605) xor estimated(607) xor estimated(637) xor estimated(639);
partial_sums(8)(374) <= estimated(349) xor estimated(351) xor estimated(381) xor estimated(383);
partial_sums(8)(375) <= estimated(861) xor estimated(863) xor estimated(893) xor estimated(895);
partial_sums(8)(376) <= estimated(61) xor estimated(63) xor estimated(125) xor estimated(127);
partial_sums(8)(377) <= estimated(573) xor estimated(575) xor estimated(637) xor estimated(639);
partial_sums(8)(378) <= estimated(317) xor estimated(319) xor estimated(381) xor estimated(383);
partial_sums(8)(379) <= estimated(829) xor estimated(831) xor estimated(893) xor estimated(895);
partial_sums(8)(380) <= estimated(125) xor estimated(127);
partial_sums(8)(381) <= estimated(637) xor estimated(639);
partial_sums(8)(382) <= estimated(381) xor estimated(383);
partial_sums(8)(383) <= estimated(893) xor estimated(895);
partial_sums(8)(384) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(385) <= estimated(515) xor estimated(519) xor estimated(523) xor estimated(527) xor estimated(531) xor estimated(535) xor estimated(539) xor estimated(543) xor estimated(547) xor estimated(551) xor estimated(555) xor estimated(559) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(579) xor estimated(583) xor estimated(587) xor estimated(591) xor estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(386) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(387) <= estimated(771) xor estimated(775) xor estimated(779) xor estimated(783) xor estimated(787) xor estimated(791) xor estimated(795) xor estimated(799) xor estimated(803) xor estimated(807) xor estimated(811) xor estimated(815) xor estimated(819) xor estimated(823) xor estimated(827) xor estimated(831) xor estimated(835) xor estimated(839) xor estimated(843) xor estimated(847) xor estimated(851) xor estimated(855) xor estimated(859) xor estimated(863) xor estimated(867) xor estimated(871) xor estimated(875) xor estimated(879) xor estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(388) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(389) <= estimated(579) xor estimated(583) xor estimated(587) xor estimated(591) xor estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(390) <= estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(391) <= estimated(835) xor estimated(839) xor estimated(843) xor estimated(847) xor estimated(851) xor estimated(855) xor estimated(859) xor estimated(863) xor estimated(867) xor estimated(871) xor estimated(875) xor estimated(879) xor estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(392) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(393) <= estimated(547) xor estimated(551) xor estimated(555) xor estimated(559) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(394) <= estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(395) <= estimated(803) xor estimated(807) xor estimated(811) xor estimated(815) xor estimated(819) xor estimated(823) xor estimated(827) xor estimated(831) xor estimated(867) xor estimated(871) xor estimated(875) xor estimated(879) xor estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(396) <= estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(397) <= estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(398) <= estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(399) <= estimated(867) xor estimated(871) xor estimated(875) xor estimated(879) xor estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(400) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(401) <= estimated(531) xor estimated(535) xor estimated(539) xor estimated(543) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(402) <= estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(403) <= estimated(787) xor estimated(791) xor estimated(795) xor estimated(799) xor estimated(819) xor estimated(823) xor estimated(827) xor estimated(831) xor estimated(851) xor estimated(855) xor estimated(859) xor estimated(863) xor estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(404) <= estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(405) <= estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(406) <= estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(407) <= estimated(851) xor estimated(855) xor estimated(859) xor estimated(863) xor estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(408) <= estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(409) <= estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(410) <= estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(411) <= estimated(819) xor estimated(823) xor estimated(827) xor estimated(831) xor estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(412) <= estimated(115) xor estimated(119) xor estimated(123) xor estimated(127);
partial_sums(8)(413) <= estimated(627) xor estimated(631) xor estimated(635) xor estimated(639);
partial_sums(8)(414) <= estimated(371) xor estimated(375) xor estimated(379) xor estimated(383);
partial_sums(8)(415) <= estimated(883) xor estimated(887) xor estimated(891) xor estimated(895);
partial_sums(8)(416) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31) xor estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(417) <= estimated(523) xor estimated(527) xor estimated(539) xor estimated(543) xor estimated(555) xor estimated(559) xor estimated(571) xor estimated(575) xor estimated(587) xor estimated(591) xor estimated(603) xor estimated(607) xor estimated(619) xor estimated(623) xor estimated(635) xor estimated(639);
partial_sums(8)(418) <= estimated(267) xor estimated(271) xor estimated(283) xor estimated(287) xor estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(419) <= estimated(779) xor estimated(783) xor estimated(795) xor estimated(799) xor estimated(811) xor estimated(815) xor estimated(827) xor estimated(831) xor estimated(843) xor estimated(847) xor estimated(859) xor estimated(863) xor estimated(875) xor estimated(879) xor estimated(891) xor estimated(895);
partial_sums(8)(420) <= estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(421) <= estimated(587) xor estimated(591) xor estimated(603) xor estimated(607) xor estimated(619) xor estimated(623) xor estimated(635) xor estimated(639);
partial_sums(8)(422) <= estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(423) <= estimated(843) xor estimated(847) xor estimated(859) xor estimated(863) xor estimated(875) xor estimated(879) xor estimated(891) xor estimated(895);
partial_sums(8)(424) <= estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(425) <= estimated(555) xor estimated(559) xor estimated(571) xor estimated(575) xor estimated(619) xor estimated(623) xor estimated(635) xor estimated(639);
partial_sums(8)(426) <= estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(427) <= estimated(811) xor estimated(815) xor estimated(827) xor estimated(831) xor estimated(875) xor estimated(879) xor estimated(891) xor estimated(895);
partial_sums(8)(428) <= estimated(107) xor estimated(111) xor estimated(123) xor estimated(127);
partial_sums(8)(429) <= estimated(619) xor estimated(623) xor estimated(635) xor estimated(639);
partial_sums(8)(430) <= estimated(363) xor estimated(367) xor estimated(379) xor estimated(383);
partial_sums(8)(431) <= estimated(875) xor estimated(879) xor estimated(891) xor estimated(895);
partial_sums(8)(432) <= estimated(27) xor estimated(31) xor estimated(59) xor estimated(63) xor estimated(91) xor estimated(95) xor estimated(123) xor estimated(127);
partial_sums(8)(433) <= estimated(539) xor estimated(543) xor estimated(571) xor estimated(575) xor estimated(603) xor estimated(607) xor estimated(635) xor estimated(639);
partial_sums(8)(434) <= estimated(283) xor estimated(287) xor estimated(315) xor estimated(319) xor estimated(347) xor estimated(351) xor estimated(379) xor estimated(383);
partial_sums(8)(435) <= estimated(795) xor estimated(799) xor estimated(827) xor estimated(831) xor estimated(859) xor estimated(863) xor estimated(891) xor estimated(895);
partial_sums(8)(436) <= estimated(91) xor estimated(95) xor estimated(123) xor estimated(127);
partial_sums(8)(437) <= estimated(603) xor estimated(607) xor estimated(635) xor estimated(639);
partial_sums(8)(438) <= estimated(347) xor estimated(351) xor estimated(379) xor estimated(383);
partial_sums(8)(439) <= estimated(859) xor estimated(863) xor estimated(891) xor estimated(895);
partial_sums(8)(440) <= estimated(59) xor estimated(63) xor estimated(123) xor estimated(127);
partial_sums(8)(441) <= estimated(571) xor estimated(575) xor estimated(635) xor estimated(639);
partial_sums(8)(442) <= estimated(315) xor estimated(319) xor estimated(379) xor estimated(383);
partial_sums(8)(443) <= estimated(827) xor estimated(831) xor estimated(891) xor estimated(895);
partial_sums(8)(444) <= estimated(123) xor estimated(127);
partial_sums(8)(445) <= estimated(635) xor estimated(639);
partial_sums(8)(446) <= estimated(379) xor estimated(383);
partial_sums(8)(447) <= estimated(891) xor estimated(895);
partial_sums(8)(448) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31) xor estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(449) <= estimated(519) xor estimated(527) xor estimated(535) xor estimated(543) xor estimated(551) xor estimated(559) xor estimated(567) xor estimated(575) xor estimated(583) xor estimated(591) xor estimated(599) xor estimated(607) xor estimated(615) xor estimated(623) xor estimated(631) xor estimated(639);
partial_sums(8)(450) <= estimated(263) xor estimated(271) xor estimated(279) xor estimated(287) xor estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(451) <= estimated(775) xor estimated(783) xor estimated(791) xor estimated(799) xor estimated(807) xor estimated(815) xor estimated(823) xor estimated(831) xor estimated(839) xor estimated(847) xor estimated(855) xor estimated(863) xor estimated(871) xor estimated(879) xor estimated(887) xor estimated(895);
partial_sums(8)(452) <= estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(453) <= estimated(583) xor estimated(591) xor estimated(599) xor estimated(607) xor estimated(615) xor estimated(623) xor estimated(631) xor estimated(639);
partial_sums(8)(454) <= estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(455) <= estimated(839) xor estimated(847) xor estimated(855) xor estimated(863) xor estimated(871) xor estimated(879) xor estimated(887) xor estimated(895);
partial_sums(8)(456) <= estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(457) <= estimated(551) xor estimated(559) xor estimated(567) xor estimated(575) xor estimated(615) xor estimated(623) xor estimated(631) xor estimated(639);
partial_sums(8)(458) <= estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(459) <= estimated(807) xor estimated(815) xor estimated(823) xor estimated(831) xor estimated(871) xor estimated(879) xor estimated(887) xor estimated(895);
partial_sums(8)(460) <= estimated(103) xor estimated(111) xor estimated(119) xor estimated(127);
partial_sums(8)(461) <= estimated(615) xor estimated(623) xor estimated(631) xor estimated(639);
partial_sums(8)(462) <= estimated(359) xor estimated(367) xor estimated(375) xor estimated(383);
partial_sums(8)(463) <= estimated(871) xor estimated(879) xor estimated(887) xor estimated(895);
partial_sums(8)(464) <= estimated(23) xor estimated(31) xor estimated(55) xor estimated(63) xor estimated(87) xor estimated(95) xor estimated(119) xor estimated(127);
partial_sums(8)(465) <= estimated(535) xor estimated(543) xor estimated(567) xor estimated(575) xor estimated(599) xor estimated(607) xor estimated(631) xor estimated(639);
partial_sums(8)(466) <= estimated(279) xor estimated(287) xor estimated(311) xor estimated(319) xor estimated(343) xor estimated(351) xor estimated(375) xor estimated(383);
partial_sums(8)(467) <= estimated(791) xor estimated(799) xor estimated(823) xor estimated(831) xor estimated(855) xor estimated(863) xor estimated(887) xor estimated(895);
partial_sums(8)(468) <= estimated(87) xor estimated(95) xor estimated(119) xor estimated(127);
partial_sums(8)(469) <= estimated(599) xor estimated(607) xor estimated(631) xor estimated(639);
partial_sums(8)(470) <= estimated(343) xor estimated(351) xor estimated(375) xor estimated(383);
partial_sums(8)(471) <= estimated(855) xor estimated(863) xor estimated(887) xor estimated(895);
partial_sums(8)(472) <= estimated(55) xor estimated(63) xor estimated(119) xor estimated(127);
partial_sums(8)(473) <= estimated(567) xor estimated(575) xor estimated(631) xor estimated(639);
partial_sums(8)(474) <= estimated(311) xor estimated(319) xor estimated(375) xor estimated(383);
partial_sums(8)(475) <= estimated(823) xor estimated(831) xor estimated(887) xor estimated(895);
partial_sums(8)(476) <= estimated(119) xor estimated(127);
partial_sums(8)(477) <= estimated(631) xor estimated(639);
partial_sums(8)(478) <= estimated(375) xor estimated(383);
partial_sums(8)(479) <= estimated(887) xor estimated(895);
partial_sums(8)(480) <= estimated(15) xor estimated(31) xor estimated(47) xor estimated(63) xor estimated(79) xor estimated(95) xor estimated(111) xor estimated(127);
partial_sums(8)(481) <= estimated(527) xor estimated(543) xor estimated(559) xor estimated(575) xor estimated(591) xor estimated(607) xor estimated(623) xor estimated(639);
partial_sums(8)(482) <= estimated(271) xor estimated(287) xor estimated(303) xor estimated(319) xor estimated(335) xor estimated(351) xor estimated(367) xor estimated(383);
partial_sums(8)(483) <= estimated(783) xor estimated(799) xor estimated(815) xor estimated(831) xor estimated(847) xor estimated(863) xor estimated(879) xor estimated(895);
partial_sums(8)(484) <= estimated(79) xor estimated(95) xor estimated(111) xor estimated(127);
partial_sums(8)(485) <= estimated(591) xor estimated(607) xor estimated(623) xor estimated(639);
partial_sums(8)(486) <= estimated(335) xor estimated(351) xor estimated(367) xor estimated(383);
partial_sums(8)(487) <= estimated(847) xor estimated(863) xor estimated(879) xor estimated(895);
partial_sums(8)(488) <= estimated(47) xor estimated(63) xor estimated(111) xor estimated(127);
partial_sums(8)(489) <= estimated(559) xor estimated(575) xor estimated(623) xor estimated(639);
partial_sums(8)(490) <= estimated(303) xor estimated(319) xor estimated(367) xor estimated(383);
partial_sums(8)(491) <= estimated(815) xor estimated(831) xor estimated(879) xor estimated(895);
partial_sums(8)(492) <= estimated(111) xor estimated(127);
partial_sums(8)(493) <= estimated(623) xor estimated(639);
partial_sums(8)(494) <= estimated(367) xor estimated(383);
partial_sums(8)(495) <= estimated(879) xor estimated(895);
partial_sums(8)(496) <= estimated(31) xor estimated(63) xor estimated(95) xor estimated(127);
partial_sums(8)(497) <= estimated(543) xor estimated(575) xor estimated(607) xor estimated(639);
partial_sums(8)(498) <= estimated(287) xor estimated(319) xor estimated(351) xor estimated(383);
partial_sums(8)(499) <= estimated(799) xor estimated(831) xor estimated(863) xor estimated(895);
partial_sums(8)(500) <= estimated(95) xor estimated(127);
partial_sums(8)(501) <= estimated(607) xor estimated(639);
partial_sums(8)(502) <= estimated(351) xor estimated(383);
partial_sums(8)(503) <= estimated(863) xor estimated(895);
partial_sums(8)(504) <= estimated(63) xor estimated(127);
partial_sums(8)(505) <= estimated(575) xor estimated(639);
partial_sums(8)(506) <= estimated(319) xor estimated(383);
partial_sums(8)(507) <= estimated(831) xor estimated(895);
partial_sums(8)(508) <= estimated(127);
partial_sums(8)(509) <= estimated(639);
partial_sums(8)(510) <= estimated(383);
partial_sums(8)(511) <= estimated(895);
partial_sums(9)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(1) <= estimated(512) xor estimated(513) xor estimated(514) xor estimated(515) xor estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(576) xor estimated(577) xor estimated(578) xor estimated(579) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(640) xor estimated(641) xor estimated(642) xor estimated(643) xor estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(704) xor estimated(705) xor estimated(706) xor estimated(707) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(2) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(3) <= estimated(640) xor estimated(641) xor estimated(642) xor estimated(643) xor estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(704) xor estimated(705) xor estimated(706) xor estimated(707) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(4) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(5) <= estimated(576) xor estimated(577) xor estimated(578) xor estimated(579) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(704) xor estimated(705) xor estimated(706) xor estimated(707) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(6) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(7) <= estimated(704) xor estimated(705) xor estimated(706) xor estimated(707) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(8) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(9) <= estimated(544) xor estimated(545) xor estimated(546) xor estimated(547) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(10) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(11) <= estimated(672) xor estimated(673) xor estimated(674) xor estimated(675) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(12) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(13) <= estimated(608) xor estimated(609) xor estimated(610) xor estimated(611) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(14) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(15) <= estimated(736) xor estimated(737) xor estimated(738) xor estimated(739) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(16) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(17) <= estimated(528) xor estimated(529) xor estimated(530) xor estimated(531) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(18) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(19) <= estimated(656) xor estimated(657) xor estimated(658) xor estimated(659) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(20) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(21) <= estimated(592) xor estimated(593) xor estimated(594) xor estimated(595) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(22) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(23) <= estimated(720) xor estimated(721) xor estimated(722) xor estimated(723) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(24) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(25) <= estimated(560) xor estimated(561) xor estimated(562) xor estimated(563) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(26) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(27) <= estimated(688) xor estimated(689) xor estimated(690) xor estimated(691) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(28) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(29) <= estimated(624) xor estimated(625) xor estimated(626) xor estimated(627) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(30) <= estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(31) <= estimated(752) xor estimated(753) xor estimated(754) xor estimated(755) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(32) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(33) <= estimated(520) xor estimated(521) xor estimated(522) xor estimated(523) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(34) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(35) <= estimated(648) xor estimated(649) xor estimated(650) xor estimated(651) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(36) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(37) <= estimated(584) xor estimated(585) xor estimated(586) xor estimated(587) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(38) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(39) <= estimated(712) xor estimated(713) xor estimated(714) xor estimated(715) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(40) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(41) <= estimated(552) xor estimated(553) xor estimated(554) xor estimated(555) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(42) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(43) <= estimated(680) xor estimated(681) xor estimated(682) xor estimated(683) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(44) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(45) <= estimated(616) xor estimated(617) xor estimated(618) xor estimated(619) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(46) <= estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(47) <= estimated(744) xor estimated(745) xor estimated(746) xor estimated(747) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(48) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(49) <= estimated(536) xor estimated(537) xor estimated(538) xor estimated(539) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(50) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(51) <= estimated(664) xor estimated(665) xor estimated(666) xor estimated(667) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(52) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(53) <= estimated(600) xor estimated(601) xor estimated(602) xor estimated(603) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(54) <= estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(55) <= estimated(728) xor estimated(729) xor estimated(730) xor estimated(731) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(56) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(57) <= estimated(568) xor estimated(569) xor estimated(570) xor estimated(571) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(58) <= estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(59) <= estimated(696) xor estimated(697) xor estimated(698) xor estimated(699) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(60) <= estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(61) <= estimated(632) xor estimated(633) xor estimated(634) xor estimated(635) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(62) <= estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(63) <= estimated(760) xor estimated(761) xor estimated(762) xor estimated(763) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(64) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(65) <= estimated(516) xor estimated(517) xor estimated(518) xor estimated(519) xor estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(66) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(67) <= estimated(644) xor estimated(645) xor estimated(646) xor estimated(647) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(68) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(69) <= estimated(580) xor estimated(581) xor estimated(582) xor estimated(583) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(70) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(71) <= estimated(708) xor estimated(709) xor estimated(710) xor estimated(711) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(72) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(73) <= estimated(548) xor estimated(549) xor estimated(550) xor estimated(551) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(74) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(75) <= estimated(676) xor estimated(677) xor estimated(678) xor estimated(679) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(76) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(77) <= estimated(612) xor estimated(613) xor estimated(614) xor estimated(615) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(78) <= estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(79) <= estimated(740) xor estimated(741) xor estimated(742) xor estimated(743) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(80) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(81) <= estimated(532) xor estimated(533) xor estimated(534) xor estimated(535) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(82) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(83) <= estimated(660) xor estimated(661) xor estimated(662) xor estimated(663) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(84) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(85) <= estimated(596) xor estimated(597) xor estimated(598) xor estimated(599) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(86) <= estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(87) <= estimated(724) xor estimated(725) xor estimated(726) xor estimated(727) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(88) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(89) <= estimated(564) xor estimated(565) xor estimated(566) xor estimated(567) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(90) <= estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(91) <= estimated(692) xor estimated(693) xor estimated(694) xor estimated(695) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(92) <= estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(93) <= estimated(628) xor estimated(629) xor estimated(630) xor estimated(631) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(94) <= estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(95) <= estimated(756) xor estimated(757) xor estimated(758) xor estimated(759) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(96) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(97) <= estimated(524) xor estimated(525) xor estimated(526) xor estimated(527) xor estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(98) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(99) <= estimated(652) xor estimated(653) xor estimated(654) xor estimated(655) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(100) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(101) <= estimated(588) xor estimated(589) xor estimated(590) xor estimated(591) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(102) <= estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(103) <= estimated(716) xor estimated(717) xor estimated(718) xor estimated(719) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(104) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(105) <= estimated(556) xor estimated(557) xor estimated(558) xor estimated(559) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(106) <= estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(107) <= estimated(684) xor estimated(685) xor estimated(686) xor estimated(687) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(108) <= estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(109) <= estimated(620) xor estimated(621) xor estimated(622) xor estimated(623) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(110) <= estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(111) <= estimated(748) xor estimated(749) xor estimated(750) xor estimated(751) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(112) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(113) <= estimated(540) xor estimated(541) xor estimated(542) xor estimated(543) xor estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(114) <= estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(115) <= estimated(668) xor estimated(669) xor estimated(670) xor estimated(671) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(116) <= estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(117) <= estimated(604) xor estimated(605) xor estimated(606) xor estimated(607) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(118) <= estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(119) <= estimated(732) xor estimated(733) xor estimated(734) xor estimated(735) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(120) <= estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(121) <= estimated(572) xor estimated(573) xor estimated(574) xor estimated(575) xor estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(122) <= estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(123) <= estimated(700) xor estimated(701) xor estimated(702) xor estimated(703) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(124) <= estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(125) <= estimated(636) xor estimated(637) xor estimated(638) xor estimated(639) xor estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(126) <= estimated(252) xor estimated(253) xor estimated(254) xor estimated(255);
partial_sums(9)(127) <= estimated(764) xor estimated(765) xor estimated(766) xor estimated(767);
partial_sums(9)(128) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(129) <= estimated(514) xor estimated(515) xor estimated(518) xor estimated(519) xor estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(546) xor estimated(547) xor estimated(550) xor estimated(551) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(578) xor estimated(579) xor estimated(582) xor estimated(583) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(642) xor estimated(643) xor estimated(646) xor estimated(647) xor estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(674) xor estimated(675) xor estimated(678) xor estimated(679) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(706) xor estimated(707) xor estimated(710) xor estimated(711) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(130) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(131) <= estimated(642) xor estimated(643) xor estimated(646) xor estimated(647) xor estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(674) xor estimated(675) xor estimated(678) xor estimated(679) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(706) xor estimated(707) xor estimated(710) xor estimated(711) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(132) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(133) <= estimated(578) xor estimated(579) xor estimated(582) xor estimated(583) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(706) xor estimated(707) xor estimated(710) xor estimated(711) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(134) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(135) <= estimated(706) xor estimated(707) xor estimated(710) xor estimated(711) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(136) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(137) <= estimated(546) xor estimated(547) xor estimated(550) xor estimated(551) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(674) xor estimated(675) xor estimated(678) xor estimated(679) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(138) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(139) <= estimated(674) xor estimated(675) xor estimated(678) xor estimated(679) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(140) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(141) <= estimated(610) xor estimated(611) xor estimated(614) xor estimated(615) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(142) <= estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(143) <= estimated(738) xor estimated(739) xor estimated(742) xor estimated(743) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(144) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(145) <= estimated(530) xor estimated(531) xor estimated(534) xor estimated(535) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(146) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(147) <= estimated(658) xor estimated(659) xor estimated(662) xor estimated(663) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(148) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(149) <= estimated(594) xor estimated(595) xor estimated(598) xor estimated(599) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(150) <= estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(151) <= estimated(722) xor estimated(723) xor estimated(726) xor estimated(727) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(152) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(153) <= estimated(562) xor estimated(563) xor estimated(566) xor estimated(567) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(154) <= estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(155) <= estimated(690) xor estimated(691) xor estimated(694) xor estimated(695) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(156) <= estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(157) <= estimated(626) xor estimated(627) xor estimated(630) xor estimated(631) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(158) <= estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(159) <= estimated(754) xor estimated(755) xor estimated(758) xor estimated(759) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(160) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(161) <= estimated(522) xor estimated(523) xor estimated(526) xor estimated(527) xor estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(162) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(163) <= estimated(650) xor estimated(651) xor estimated(654) xor estimated(655) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(164) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(165) <= estimated(586) xor estimated(587) xor estimated(590) xor estimated(591) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(166) <= estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(167) <= estimated(714) xor estimated(715) xor estimated(718) xor estimated(719) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(168) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(169) <= estimated(554) xor estimated(555) xor estimated(558) xor estimated(559) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(170) <= estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(171) <= estimated(682) xor estimated(683) xor estimated(686) xor estimated(687) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(172) <= estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(173) <= estimated(618) xor estimated(619) xor estimated(622) xor estimated(623) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(174) <= estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(175) <= estimated(746) xor estimated(747) xor estimated(750) xor estimated(751) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(176) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(177) <= estimated(538) xor estimated(539) xor estimated(542) xor estimated(543) xor estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(178) <= estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(179) <= estimated(666) xor estimated(667) xor estimated(670) xor estimated(671) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(180) <= estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(181) <= estimated(602) xor estimated(603) xor estimated(606) xor estimated(607) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(182) <= estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(183) <= estimated(730) xor estimated(731) xor estimated(734) xor estimated(735) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(184) <= estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(185) <= estimated(570) xor estimated(571) xor estimated(574) xor estimated(575) xor estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(186) <= estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(187) <= estimated(698) xor estimated(699) xor estimated(702) xor estimated(703) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(188) <= estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(189) <= estimated(634) xor estimated(635) xor estimated(638) xor estimated(639) xor estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(190) <= estimated(250) xor estimated(251) xor estimated(254) xor estimated(255);
partial_sums(9)(191) <= estimated(762) xor estimated(763) xor estimated(766) xor estimated(767);
partial_sums(9)(192) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(193) <= estimated(518) xor estimated(519) xor estimated(526) xor estimated(527) xor estimated(534) xor estimated(535) xor estimated(542) xor estimated(543) xor estimated(550) xor estimated(551) xor estimated(558) xor estimated(559) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(582) xor estimated(583) xor estimated(590) xor estimated(591) xor estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(646) xor estimated(647) xor estimated(654) xor estimated(655) xor estimated(662) xor estimated(663) xor estimated(670) xor estimated(671) xor estimated(678) xor estimated(679) xor estimated(686) xor estimated(687) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(710) xor estimated(711) xor estimated(718) xor estimated(719) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(194) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(195) <= estimated(646) xor estimated(647) xor estimated(654) xor estimated(655) xor estimated(662) xor estimated(663) xor estimated(670) xor estimated(671) xor estimated(678) xor estimated(679) xor estimated(686) xor estimated(687) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(710) xor estimated(711) xor estimated(718) xor estimated(719) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(196) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(197) <= estimated(582) xor estimated(583) xor estimated(590) xor estimated(591) xor estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(710) xor estimated(711) xor estimated(718) xor estimated(719) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(198) <= estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(199) <= estimated(710) xor estimated(711) xor estimated(718) xor estimated(719) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(200) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(201) <= estimated(550) xor estimated(551) xor estimated(558) xor estimated(559) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(678) xor estimated(679) xor estimated(686) xor estimated(687) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(202) <= estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(203) <= estimated(678) xor estimated(679) xor estimated(686) xor estimated(687) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(204) <= estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(205) <= estimated(614) xor estimated(615) xor estimated(622) xor estimated(623) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(206) <= estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(207) <= estimated(742) xor estimated(743) xor estimated(750) xor estimated(751) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(208) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(209) <= estimated(534) xor estimated(535) xor estimated(542) xor estimated(543) xor estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(662) xor estimated(663) xor estimated(670) xor estimated(671) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(210) <= estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(211) <= estimated(662) xor estimated(663) xor estimated(670) xor estimated(671) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(212) <= estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(213) <= estimated(598) xor estimated(599) xor estimated(606) xor estimated(607) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(214) <= estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(215) <= estimated(726) xor estimated(727) xor estimated(734) xor estimated(735) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(216) <= estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(217) <= estimated(566) xor estimated(567) xor estimated(574) xor estimated(575) xor estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(218) <= estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(219) <= estimated(694) xor estimated(695) xor estimated(702) xor estimated(703) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(220) <= estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(221) <= estimated(630) xor estimated(631) xor estimated(638) xor estimated(639) xor estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(222) <= estimated(246) xor estimated(247) xor estimated(254) xor estimated(255);
partial_sums(9)(223) <= estimated(758) xor estimated(759) xor estimated(766) xor estimated(767);
partial_sums(9)(224) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31) xor estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(225) <= estimated(526) xor estimated(527) xor estimated(542) xor estimated(543) xor estimated(558) xor estimated(559) xor estimated(574) xor estimated(575) xor estimated(590) xor estimated(591) xor estimated(606) xor estimated(607) xor estimated(622) xor estimated(623) xor estimated(638) xor estimated(639) xor estimated(654) xor estimated(655) xor estimated(670) xor estimated(671) xor estimated(686) xor estimated(687) xor estimated(702) xor estimated(703) xor estimated(718) xor estimated(719) xor estimated(734) xor estimated(735) xor estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(226) <= estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(227) <= estimated(654) xor estimated(655) xor estimated(670) xor estimated(671) xor estimated(686) xor estimated(687) xor estimated(702) xor estimated(703) xor estimated(718) xor estimated(719) xor estimated(734) xor estimated(735) xor estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(228) <= estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(229) <= estimated(590) xor estimated(591) xor estimated(606) xor estimated(607) xor estimated(622) xor estimated(623) xor estimated(638) xor estimated(639) xor estimated(718) xor estimated(719) xor estimated(734) xor estimated(735) xor estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(230) <= estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(231) <= estimated(718) xor estimated(719) xor estimated(734) xor estimated(735) xor estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(232) <= estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(233) <= estimated(558) xor estimated(559) xor estimated(574) xor estimated(575) xor estimated(622) xor estimated(623) xor estimated(638) xor estimated(639) xor estimated(686) xor estimated(687) xor estimated(702) xor estimated(703) xor estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(234) <= estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(235) <= estimated(686) xor estimated(687) xor estimated(702) xor estimated(703) xor estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(236) <= estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(237) <= estimated(622) xor estimated(623) xor estimated(638) xor estimated(639) xor estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(238) <= estimated(238) xor estimated(239) xor estimated(254) xor estimated(255);
partial_sums(9)(239) <= estimated(750) xor estimated(751) xor estimated(766) xor estimated(767);
partial_sums(9)(240) <= estimated(30) xor estimated(31) xor estimated(62) xor estimated(63) xor estimated(94) xor estimated(95) xor estimated(126) xor estimated(127) xor estimated(158) xor estimated(159) xor estimated(190) xor estimated(191) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(241) <= estimated(542) xor estimated(543) xor estimated(574) xor estimated(575) xor estimated(606) xor estimated(607) xor estimated(638) xor estimated(639) xor estimated(670) xor estimated(671) xor estimated(702) xor estimated(703) xor estimated(734) xor estimated(735) xor estimated(766) xor estimated(767);
partial_sums(9)(242) <= estimated(158) xor estimated(159) xor estimated(190) xor estimated(191) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(243) <= estimated(670) xor estimated(671) xor estimated(702) xor estimated(703) xor estimated(734) xor estimated(735) xor estimated(766) xor estimated(767);
partial_sums(9)(244) <= estimated(94) xor estimated(95) xor estimated(126) xor estimated(127) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(245) <= estimated(606) xor estimated(607) xor estimated(638) xor estimated(639) xor estimated(734) xor estimated(735) xor estimated(766) xor estimated(767);
partial_sums(9)(246) <= estimated(222) xor estimated(223) xor estimated(254) xor estimated(255);
partial_sums(9)(247) <= estimated(734) xor estimated(735) xor estimated(766) xor estimated(767);
partial_sums(9)(248) <= estimated(62) xor estimated(63) xor estimated(126) xor estimated(127) xor estimated(190) xor estimated(191) xor estimated(254) xor estimated(255);
partial_sums(9)(249) <= estimated(574) xor estimated(575) xor estimated(638) xor estimated(639) xor estimated(702) xor estimated(703) xor estimated(766) xor estimated(767);
partial_sums(9)(250) <= estimated(190) xor estimated(191) xor estimated(254) xor estimated(255);
partial_sums(9)(251) <= estimated(702) xor estimated(703) xor estimated(766) xor estimated(767);
partial_sums(9)(252) <= estimated(126) xor estimated(127) xor estimated(254) xor estimated(255);
partial_sums(9)(253) <= estimated(638) xor estimated(639) xor estimated(766) xor estimated(767);
partial_sums(9)(254) <= estimated(254) xor estimated(255);
partial_sums(9)(255) <= estimated(766) xor estimated(767);
partial_sums(9)(256) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(257) <= estimated(513) xor estimated(515) xor estimated(517) xor estimated(519) xor estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(545) xor estimated(547) xor estimated(549) xor estimated(551) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(577) xor estimated(579) xor estimated(581) xor estimated(583) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(641) xor estimated(643) xor estimated(645) xor estimated(647) xor estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(673) xor estimated(675) xor estimated(677) xor estimated(679) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(705) xor estimated(707) xor estimated(709) xor estimated(711) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(258) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(259) <= estimated(641) xor estimated(643) xor estimated(645) xor estimated(647) xor estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(673) xor estimated(675) xor estimated(677) xor estimated(679) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(705) xor estimated(707) xor estimated(709) xor estimated(711) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(260) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(261) <= estimated(577) xor estimated(579) xor estimated(581) xor estimated(583) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(705) xor estimated(707) xor estimated(709) xor estimated(711) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(262) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(263) <= estimated(705) xor estimated(707) xor estimated(709) xor estimated(711) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(264) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(265) <= estimated(545) xor estimated(547) xor estimated(549) xor estimated(551) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(673) xor estimated(675) xor estimated(677) xor estimated(679) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(266) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(267) <= estimated(673) xor estimated(675) xor estimated(677) xor estimated(679) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(268) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(269) <= estimated(609) xor estimated(611) xor estimated(613) xor estimated(615) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(270) <= estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(271) <= estimated(737) xor estimated(739) xor estimated(741) xor estimated(743) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(272) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(273) <= estimated(529) xor estimated(531) xor estimated(533) xor estimated(535) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(274) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(275) <= estimated(657) xor estimated(659) xor estimated(661) xor estimated(663) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(276) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(277) <= estimated(593) xor estimated(595) xor estimated(597) xor estimated(599) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(278) <= estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(279) <= estimated(721) xor estimated(723) xor estimated(725) xor estimated(727) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(280) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(281) <= estimated(561) xor estimated(563) xor estimated(565) xor estimated(567) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(282) <= estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(283) <= estimated(689) xor estimated(691) xor estimated(693) xor estimated(695) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(284) <= estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(285) <= estimated(625) xor estimated(627) xor estimated(629) xor estimated(631) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(286) <= estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(287) <= estimated(753) xor estimated(755) xor estimated(757) xor estimated(759) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(288) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(289) <= estimated(521) xor estimated(523) xor estimated(525) xor estimated(527) xor estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(290) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(291) <= estimated(649) xor estimated(651) xor estimated(653) xor estimated(655) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(292) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(293) <= estimated(585) xor estimated(587) xor estimated(589) xor estimated(591) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(294) <= estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(295) <= estimated(713) xor estimated(715) xor estimated(717) xor estimated(719) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(296) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(297) <= estimated(553) xor estimated(555) xor estimated(557) xor estimated(559) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(298) <= estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(299) <= estimated(681) xor estimated(683) xor estimated(685) xor estimated(687) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(300) <= estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(301) <= estimated(617) xor estimated(619) xor estimated(621) xor estimated(623) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(302) <= estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(303) <= estimated(745) xor estimated(747) xor estimated(749) xor estimated(751) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(304) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(305) <= estimated(537) xor estimated(539) xor estimated(541) xor estimated(543) xor estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(306) <= estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(307) <= estimated(665) xor estimated(667) xor estimated(669) xor estimated(671) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(308) <= estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(309) <= estimated(601) xor estimated(603) xor estimated(605) xor estimated(607) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(310) <= estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(311) <= estimated(729) xor estimated(731) xor estimated(733) xor estimated(735) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(312) <= estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(313) <= estimated(569) xor estimated(571) xor estimated(573) xor estimated(575) xor estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(314) <= estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(315) <= estimated(697) xor estimated(699) xor estimated(701) xor estimated(703) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(316) <= estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(317) <= estimated(633) xor estimated(635) xor estimated(637) xor estimated(639) xor estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(318) <= estimated(249) xor estimated(251) xor estimated(253) xor estimated(255);
partial_sums(9)(319) <= estimated(761) xor estimated(763) xor estimated(765) xor estimated(767);
partial_sums(9)(320) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(321) <= estimated(517) xor estimated(519) xor estimated(525) xor estimated(527) xor estimated(533) xor estimated(535) xor estimated(541) xor estimated(543) xor estimated(549) xor estimated(551) xor estimated(557) xor estimated(559) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(581) xor estimated(583) xor estimated(589) xor estimated(591) xor estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(645) xor estimated(647) xor estimated(653) xor estimated(655) xor estimated(661) xor estimated(663) xor estimated(669) xor estimated(671) xor estimated(677) xor estimated(679) xor estimated(685) xor estimated(687) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(709) xor estimated(711) xor estimated(717) xor estimated(719) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(322) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(323) <= estimated(645) xor estimated(647) xor estimated(653) xor estimated(655) xor estimated(661) xor estimated(663) xor estimated(669) xor estimated(671) xor estimated(677) xor estimated(679) xor estimated(685) xor estimated(687) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(709) xor estimated(711) xor estimated(717) xor estimated(719) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(324) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(325) <= estimated(581) xor estimated(583) xor estimated(589) xor estimated(591) xor estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(709) xor estimated(711) xor estimated(717) xor estimated(719) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(326) <= estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(327) <= estimated(709) xor estimated(711) xor estimated(717) xor estimated(719) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(328) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(329) <= estimated(549) xor estimated(551) xor estimated(557) xor estimated(559) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(677) xor estimated(679) xor estimated(685) xor estimated(687) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(330) <= estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(331) <= estimated(677) xor estimated(679) xor estimated(685) xor estimated(687) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(332) <= estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(333) <= estimated(613) xor estimated(615) xor estimated(621) xor estimated(623) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(334) <= estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(335) <= estimated(741) xor estimated(743) xor estimated(749) xor estimated(751) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(336) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(337) <= estimated(533) xor estimated(535) xor estimated(541) xor estimated(543) xor estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(661) xor estimated(663) xor estimated(669) xor estimated(671) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(338) <= estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(339) <= estimated(661) xor estimated(663) xor estimated(669) xor estimated(671) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(340) <= estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(341) <= estimated(597) xor estimated(599) xor estimated(605) xor estimated(607) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(342) <= estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(343) <= estimated(725) xor estimated(727) xor estimated(733) xor estimated(735) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(344) <= estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(345) <= estimated(565) xor estimated(567) xor estimated(573) xor estimated(575) xor estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(346) <= estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(347) <= estimated(693) xor estimated(695) xor estimated(701) xor estimated(703) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(348) <= estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(349) <= estimated(629) xor estimated(631) xor estimated(637) xor estimated(639) xor estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(350) <= estimated(245) xor estimated(247) xor estimated(253) xor estimated(255);
partial_sums(9)(351) <= estimated(757) xor estimated(759) xor estimated(765) xor estimated(767);
partial_sums(9)(352) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31) xor estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(353) <= estimated(525) xor estimated(527) xor estimated(541) xor estimated(543) xor estimated(557) xor estimated(559) xor estimated(573) xor estimated(575) xor estimated(589) xor estimated(591) xor estimated(605) xor estimated(607) xor estimated(621) xor estimated(623) xor estimated(637) xor estimated(639) xor estimated(653) xor estimated(655) xor estimated(669) xor estimated(671) xor estimated(685) xor estimated(687) xor estimated(701) xor estimated(703) xor estimated(717) xor estimated(719) xor estimated(733) xor estimated(735) xor estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(354) <= estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(355) <= estimated(653) xor estimated(655) xor estimated(669) xor estimated(671) xor estimated(685) xor estimated(687) xor estimated(701) xor estimated(703) xor estimated(717) xor estimated(719) xor estimated(733) xor estimated(735) xor estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(356) <= estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(357) <= estimated(589) xor estimated(591) xor estimated(605) xor estimated(607) xor estimated(621) xor estimated(623) xor estimated(637) xor estimated(639) xor estimated(717) xor estimated(719) xor estimated(733) xor estimated(735) xor estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(358) <= estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(359) <= estimated(717) xor estimated(719) xor estimated(733) xor estimated(735) xor estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(360) <= estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(361) <= estimated(557) xor estimated(559) xor estimated(573) xor estimated(575) xor estimated(621) xor estimated(623) xor estimated(637) xor estimated(639) xor estimated(685) xor estimated(687) xor estimated(701) xor estimated(703) xor estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(362) <= estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(363) <= estimated(685) xor estimated(687) xor estimated(701) xor estimated(703) xor estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(364) <= estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(365) <= estimated(621) xor estimated(623) xor estimated(637) xor estimated(639) xor estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(366) <= estimated(237) xor estimated(239) xor estimated(253) xor estimated(255);
partial_sums(9)(367) <= estimated(749) xor estimated(751) xor estimated(765) xor estimated(767);
partial_sums(9)(368) <= estimated(29) xor estimated(31) xor estimated(61) xor estimated(63) xor estimated(93) xor estimated(95) xor estimated(125) xor estimated(127) xor estimated(157) xor estimated(159) xor estimated(189) xor estimated(191) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(369) <= estimated(541) xor estimated(543) xor estimated(573) xor estimated(575) xor estimated(605) xor estimated(607) xor estimated(637) xor estimated(639) xor estimated(669) xor estimated(671) xor estimated(701) xor estimated(703) xor estimated(733) xor estimated(735) xor estimated(765) xor estimated(767);
partial_sums(9)(370) <= estimated(157) xor estimated(159) xor estimated(189) xor estimated(191) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(371) <= estimated(669) xor estimated(671) xor estimated(701) xor estimated(703) xor estimated(733) xor estimated(735) xor estimated(765) xor estimated(767);
partial_sums(9)(372) <= estimated(93) xor estimated(95) xor estimated(125) xor estimated(127) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(373) <= estimated(605) xor estimated(607) xor estimated(637) xor estimated(639) xor estimated(733) xor estimated(735) xor estimated(765) xor estimated(767);
partial_sums(9)(374) <= estimated(221) xor estimated(223) xor estimated(253) xor estimated(255);
partial_sums(9)(375) <= estimated(733) xor estimated(735) xor estimated(765) xor estimated(767);
partial_sums(9)(376) <= estimated(61) xor estimated(63) xor estimated(125) xor estimated(127) xor estimated(189) xor estimated(191) xor estimated(253) xor estimated(255);
partial_sums(9)(377) <= estimated(573) xor estimated(575) xor estimated(637) xor estimated(639) xor estimated(701) xor estimated(703) xor estimated(765) xor estimated(767);
partial_sums(9)(378) <= estimated(189) xor estimated(191) xor estimated(253) xor estimated(255);
partial_sums(9)(379) <= estimated(701) xor estimated(703) xor estimated(765) xor estimated(767);
partial_sums(9)(380) <= estimated(125) xor estimated(127) xor estimated(253) xor estimated(255);
partial_sums(9)(381) <= estimated(637) xor estimated(639) xor estimated(765) xor estimated(767);
partial_sums(9)(382) <= estimated(253) xor estimated(255);
partial_sums(9)(383) <= estimated(765) xor estimated(767);
partial_sums(9)(384) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(385) <= estimated(515) xor estimated(519) xor estimated(523) xor estimated(527) xor estimated(531) xor estimated(535) xor estimated(539) xor estimated(543) xor estimated(547) xor estimated(551) xor estimated(555) xor estimated(559) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(579) xor estimated(583) xor estimated(587) xor estimated(591) xor estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(643) xor estimated(647) xor estimated(651) xor estimated(655) xor estimated(659) xor estimated(663) xor estimated(667) xor estimated(671) xor estimated(675) xor estimated(679) xor estimated(683) xor estimated(687) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(707) xor estimated(711) xor estimated(715) xor estimated(719) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(386) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(387) <= estimated(643) xor estimated(647) xor estimated(651) xor estimated(655) xor estimated(659) xor estimated(663) xor estimated(667) xor estimated(671) xor estimated(675) xor estimated(679) xor estimated(683) xor estimated(687) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(707) xor estimated(711) xor estimated(715) xor estimated(719) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(388) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(389) <= estimated(579) xor estimated(583) xor estimated(587) xor estimated(591) xor estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(707) xor estimated(711) xor estimated(715) xor estimated(719) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(390) <= estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(391) <= estimated(707) xor estimated(711) xor estimated(715) xor estimated(719) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(392) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(393) <= estimated(547) xor estimated(551) xor estimated(555) xor estimated(559) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(675) xor estimated(679) xor estimated(683) xor estimated(687) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(394) <= estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(395) <= estimated(675) xor estimated(679) xor estimated(683) xor estimated(687) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(396) <= estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(397) <= estimated(611) xor estimated(615) xor estimated(619) xor estimated(623) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(398) <= estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(399) <= estimated(739) xor estimated(743) xor estimated(747) xor estimated(751) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(400) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(401) <= estimated(531) xor estimated(535) xor estimated(539) xor estimated(543) xor estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(659) xor estimated(663) xor estimated(667) xor estimated(671) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(402) <= estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(403) <= estimated(659) xor estimated(663) xor estimated(667) xor estimated(671) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(404) <= estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(405) <= estimated(595) xor estimated(599) xor estimated(603) xor estimated(607) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(406) <= estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(407) <= estimated(723) xor estimated(727) xor estimated(731) xor estimated(735) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(408) <= estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(409) <= estimated(563) xor estimated(567) xor estimated(571) xor estimated(575) xor estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(410) <= estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(411) <= estimated(691) xor estimated(695) xor estimated(699) xor estimated(703) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(412) <= estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(413) <= estimated(627) xor estimated(631) xor estimated(635) xor estimated(639) xor estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(414) <= estimated(243) xor estimated(247) xor estimated(251) xor estimated(255);
partial_sums(9)(415) <= estimated(755) xor estimated(759) xor estimated(763) xor estimated(767);
partial_sums(9)(416) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31) xor estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(417) <= estimated(523) xor estimated(527) xor estimated(539) xor estimated(543) xor estimated(555) xor estimated(559) xor estimated(571) xor estimated(575) xor estimated(587) xor estimated(591) xor estimated(603) xor estimated(607) xor estimated(619) xor estimated(623) xor estimated(635) xor estimated(639) xor estimated(651) xor estimated(655) xor estimated(667) xor estimated(671) xor estimated(683) xor estimated(687) xor estimated(699) xor estimated(703) xor estimated(715) xor estimated(719) xor estimated(731) xor estimated(735) xor estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(418) <= estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(419) <= estimated(651) xor estimated(655) xor estimated(667) xor estimated(671) xor estimated(683) xor estimated(687) xor estimated(699) xor estimated(703) xor estimated(715) xor estimated(719) xor estimated(731) xor estimated(735) xor estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(420) <= estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(421) <= estimated(587) xor estimated(591) xor estimated(603) xor estimated(607) xor estimated(619) xor estimated(623) xor estimated(635) xor estimated(639) xor estimated(715) xor estimated(719) xor estimated(731) xor estimated(735) xor estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(422) <= estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(423) <= estimated(715) xor estimated(719) xor estimated(731) xor estimated(735) xor estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(424) <= estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(425) <= estimated(555) xor estimated(559) xor estimated(571) xor estimated(575) xor estimated(619) xor estimated(623) xor estimated(635) xor estimated(639) xor estimated(683) xor estimated(687) xor estimated(699) xor estimated(703) xor estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(426) <= estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(427) <= estimated(683) xor estimated(687) xor estimated(699) xor estimated(703) xor estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(428) <= estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(429) <= estimated(619) xor estimated(623) xor estimated(635) xor estimated(639) xor estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(430) <= estimated(235) xor estimated(239) xor estimated(251) xor estimated(255);
partial_sums(9)(431) <= estimated(747) xor estimated(751) xor estimated(763) xor estimated(767);
partial_sums(9)(432) <= estimated(27) xor estimated(31) xor estimated(59) xor estimated(63) xor estimated(91) xor estimated(95) xor estimated(123) xor estimated(127) xor estimated(155) xor estimated(159) xor estimated(187) xor estimated(191) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(433) <= estimated(539) xor estimated(543) xor estimated(571) xor estimated(575) xor estimated(603) xor estimated(607) xor estimated(635) xor estimated(639) xor estimated(667) xor estimated(671) xor estimated(699) xor estimated(703) xor estimated(731) xor estimated(735) xor estimated(763) xor estimated(767);
partial_sums(9)(434) <= estimated(155) xor estimated(159) xor estimated(187) xor estimated(191) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(435) <= estimated(667) xor estimated(671) xor estimated(699) xor estimated(703) xor estimated(731) xor estimated(735) xor estimated(763) xor estimated(767);
partial_sums(9)(436) <= estimated(91) xor estimated(95) xor estimated(123) xor estimated(127) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(437) <= estimated(603) xor estimated(607) xor estimated(635) xor estimated(639) xor estimated(731) xor estimated(735) xor estimated(763) xor estimated(767);
partial_sums(9)(438) <= estimated(219) xor estimated(223) xor estimated(251) xor estimated(255);
partial_sums(9)(439) <= estimated(731) xor estimated(735) xor estimated(763) xor estimated(767);
partial_sums(9)(440) <= estimated(59) xor estimated(63) xor estimated(123) xor estimated(127) xor estimated(187) xor estimated(191) xor estimated(251) xor estimated(255);
partial_sums(9)(441) <= estimated(571) xor estimated(575) xor estimated(635) xor estimated(639) xor estimated(699) xor estimated(703) xor estimated(763) xor estimated(767);
partial_sums(9)(442) <= estimated(187) xor estimated(191) xor estimated(251) xor estimated(255);
partial_sums(9)(443) <= estimated(699) xor estimated(703) xor estimated(763) xor estimated(767);
partial_sums(9)(444) <= estimated(123) xor estimated(127) xor estimated(251) xor estimated(255);
partial_sums(9)(445) <= estimated(635) xor estimated(639) xor estimated(763) xor estimated(767);
partial_sums(9)(446) <= estimated(251) xor estimated(255);
partial_sums(9)(447) <= estimated(763) xor estimated(767);
partial_sums(9)(448) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31) xor estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(449) <= estimated(519) xor estimated(527) xor estimated(535) xor estimated(543) xor estimated(551) xor estimated(559) xor estimated(567) xor estimated(575) xor estimated(583) xor estimated(591) xor estimated(599) xor estimated(607) xor estimated(615) xor estimated(623) xor estimated(631) xor estimated(639) xor estimated(647) xor estimated(655) xor estimated(663) xor estimated(671) xor estimated(679) xor estimated(687) xor estimated(695) xor estimated(703) xor estimated(711) xor estimated(719) xor estimated(727) xor estimated(735) xor estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(450) <= estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(451) <= estimated(647) xor estimated(655) xor estimated(663) xor estimated(671) xor estimated(679) xor estimated(687) xor estimated(695) xor estimated(703) xor estimated(711) xor estimated(719) xor estimated(727) xor estimated(735) xor estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(452) <= estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(453) <= estimated(583) xor estimated(591) xor estimated(599) xor estimated(607) xor estimated(615) xor estimated(623) xor estimated(631) xor estimated(639) xor estimated(711) xor estimated(719) xor estimated(727) xor estimated(735) xor estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(454) <= estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(455) <= estimated(711) xor estimated(719) xor estimated(727) xor estimated(735) xor estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(456) <= estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(457) <= estimated(551) xor estimated(559) xor estimated(567) xor estimated(575) xor estimated(615) xor estimated(623) xor estimated(631) xor estimated(639) xor estimated(679) xor estimated(687) xor estimated(695) xor estimated(703) xor estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(458) <= estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(459) <= estimated(679) xor estimated(687) xor estimated(695) xor estimated(703) xor estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(460) <= estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(461) <= estimated(615) xor estimated(623) xor estimated(631) xor estimated(639) xor estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(462) <= estimated(231) xor estimated(239) xor estimated(247) xor estimated(255);
partial_sums(9)(463) <= estimated(743) xor estimated(751) xor estimated(759) xor estimated(767);
partial_sums(9)(464) <= estimated(23) xor estimated(31) xor estimated(55) xor estimated(63) xor estimated(87) xor estimated(95) xor estimated(119) xor estimated(127) xor estimated(151) xor estimated(159) xor estimated(183) xor estimated(191) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(465) <= estimated(535) xor estimated(543) xor estimated(567) xor estimated(575) xor estimated(599) xor estimated(607) xor estimated(631) xor estimated(639) xor estimated(663) xor estimated(671) xor estimated(695) xor estimated(703) xor estimated(727) xor estimated(735) xor estimated(759) xor estimated(767);
partial_sums(9)(466) <= estimated(151) xor estimated(159) xor estimated(183) xor estimated(191) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(467) <= estimated(663) xor estimated(671) xor estimated(695) xor estimated(703) xor estimated(727) xor estimated(735) xor estimated(759) xor estimated(767);
partial_sums(9)(468) <= estimated(87) xor estimated(95) xor estimated(119) xor estimated(127) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(469) <= estimated(599) xor estimated(607) xor estimated(631) xor estimated(639) xor estimated(727) xor estimated(735) xor estimated(759) xor estimated(767);
partial_sums(9)(470) <= estimated(215) xor estimated(223) xor estimated(247) xor estimated(255);
partial_sums(9)(471) <= estimated(727) xor estimated(735) xor estimated(759) xor estimated(767);
partial_sums(9)(472) <= estimated(55) xor estimated(63) xor estimated(119) xor estimated(127) xor estimated(183) xor estimated(191) xor estimated(247) xor estimated(255);
partial_sums(9)(473) <= estimated(567) xor estimated(575) xor estimated(631) xor estimated(639) xor estimated(695) xor estimated(703) xor estimated(759) xor estimated(767);
partial_sums(9)(474) <= estimated(183) xor estimated(191) xor estimated(247) xor estimated(255);
partial_sums(9)(475) <= estimated(695) xor estimated(703) xor estimated(759) xor estimated(767);
partial_sums(9)(476) <= estimated(119) xor estimated(127) xor estimated(247) xor estimated(255);
partial_sums(9)(477) <= estimated(631) xor estimated(639) xor estimated(759) xor estimated(767);
partial_sums(9)(478) <= estimated(247) xor estimated(255);
partial_sums(9)(479) <= estimated(759) xor estimated(767);
partial_sums(9)(480) <= estimated(15) xor estimated(31) xor estimated(47) xor estimated(63) xor estimated(79) xor estimated(95) xor estimated(111) xor estimated(127) xor estimated(143) xor estimated(159) xor estimated(175) xor estimated(191) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(481) <= estimated(527) xor estimated(543) xor estimated(559) xor estimated(575) xor estimated(591) xor estimated(607) xor estimated(623) xor estimated(639) xor estimated(655) xor estimated(671) xor estimated(687) xor estimated(703) xor estimated(719) xor estimated(735) xor estimated(751) xor estimated(767);
partial_sums(9)(482) <= estimated(143) xor estimated(159) xor estimated(175) xor estimated(191) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(483) <= estimated(655) xor estimated(671) xor estimated(687) xor estimated(703) xor estimated(719) xor estimated(735) xor estimated(751) xor estimated(767);
partial_sums(9)(484) <= estimated(79) xor estimated(95) xor estimated(111) xor estimated(127) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(485) <= estimated(591) xor estimated(607) xor estimated(623) xor estimated(639) xor estimated(719) xor estimated(735) xor estimated(751) xor estimated(767);
partial_sums(9)(486) <= estimated(207) xor estimated(223) xor estimated(239) xor estimated(255);
partial_sums(9)(487) <= estimated(719) xor estimated(735) xor estimated(751) xor estimated(767);
partial_sums(9)(488) <= estimated(47) xor estimated(63) xor estimated(111) xor estimated(127) xor estimated(175) xor estimated(191) xor estimated(239) xor estimated(255);
partial_sums(9)(489) <= estimated(559) xor estimated(575) xor estimated(623) xor estimated(639) xor estimated(687) xor estimated(703) xor estimated(751) xor estimated(767);
partial_sums(9)(490) <= estimated(175) xor estimated(191) xor estimated(239) xor estimated(255);
partial_sums(9)(491) <= estimated(687) xor estimated(703) xor estimated(751) xor estimated(767);
partial_sums(9)(492) <= estimated(111) xor estimated(127) xor estimated(239) xor estimated(255);
partial_sums(9)(493) <= estimated(623) xor estimated(639) xor estimated(751) xor estimated(767);
partial_sums(9)(494) <= estimated(239) xor estimated(255);
partial_sums(9)(495) <= estimated(751) xor estimated(767);
partial_sums(9)(496) <= estimated(31) xor estimated(63) xor estimated(95) xor estimated(127) xor estimated(159) xor estimated(191) xor estimated(223) xor estimated(255);
partial_sums(9)(497) <= estimated(543) xor estimated(575) xor estimated(607) xor estimated(639) xor estimated(671) xor estimated(703) xor estimated(735) xor estimated(767);
partial_sums(9)(498) <= estimated(159) xor estimated(191) xor estimated(223) xor estimated(255);
partial_sums(9)(499) <= estimated(671) xor estimated(703) xor estimated(735) xor estimated(767);
partial_sums(9)(500) <= estimated(95) xor estimated(127) xor estimated(223) xor estimated(255);
partial_sums(9)(501) <= estimated(607) xor estimated(639) xor estimated(735) xor estimated(767);
partial_sums(9)(502) <= estimated(223) xor estimated(255);
partial_sums(9)(503) <= estimated(735) xor estimated(767);
partial_sums(9)(504) <= estimated(63) xor estimated(127) xor estimated(191) xor estimated(255);
partial_sums(9)(505) <= estimated(575) xor estimated(639) xor estimated(703) xor estimated(767);
partial_sums(9)(506) <= estimated(191) xor estimated(255);
partial_sums(9)(507) <= estimated(703) xor estimated(767);
partial_sums(9)(508) <= estimated(127) xor estimated(255);
partial_sums(9)(509) <= estimated(639) xor estimated(767);
partial_sums(9)(510) <= estimated(255);
partial_sums(9)(511) <= estimated(767);
partial_sums(10)(0) <= estimated(0) xor estimated(1) xor estimated(2) xor estimated(3) xor estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(1) <= estimated(256) xor estimated(257) xor estimated(258) xor estimated(259) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(2) <= estimated(128) xor estimated(129) xor estimated(130) xor estimated(131) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(3) <= estimated(384) xor estimated(385) xor estimated(386) xor estimated(387) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(4) <= estimated(64) xor estimated(65) xor estimated(66) xor estimated(67) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(5) <= estimated(320) xor estimated(321) xor estimated(322) xor estimated(323) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(6) <= estimated(192) xor estimated(193) xor estimated(194) xor estimated(195) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(7) <= estimated(448) xor estimated(449) xor estimated(450) xor estimated(451) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(8) <= estimated(32) xor estimated(33) xor estimated(34) xor estimated(35) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(9) <= estimated(288) xor estimated(289) xor estimated(290) xor estimated(291) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(10) <= estimated(160) xor estimated(161) xor estimated(162) xor estimated(163) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(11) <= estimated(416) xor estimated(417) xor estimated(418) xor estimated(419) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(12) <= estimated(96) xor estimated(97) xor estimated(98) xor estimated(99) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(13) <= estimated(352) xor estimated(353) xor estimated(354) xor estimated(355) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(14) <= estimated(224) xor estimated(225) xor estimated(226) xor estimated(227) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(15) <= estimated(480) xor estimated(481) xor estimated(482) xor estimated(483) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(16) <= estimated(16) xor estimated(17) xor estimated(18) xor estimated(19) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(17) <= estimated(272) xor estimated(273) xor estimated(274) xor estimated(275) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(18) <= estimated(144) xor estimated(145) xor estimated(146) xor estimated(147) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(19) <= estimated(400) xor estimated(401) xor estimated(402) xor estimated(403) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(20) <= estimated(80) xor estimated(81) xor estimated(82) xor estimated(83) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(21) <= estimated(336) xor estimated(337) xor estimated(338) xor estimated(339) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(22) <= estimated(208) xor estimated(209) xor estimated(210) xor estimated(211) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(23) <= estimated(464) xor estimated(465) xor estimated(466) xor estimated(467) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(24) <= estimated(48) xor estimated(49) xor estimated(50) xor estimated(51) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(25) <= estimated(304) xor estimated(305) xor estimated(306) xor estimated(307) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(26) <= estimated(176) xor estimated(177) xor estimated(178) xor estimated(179) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(27) <= estimated(432) xor estimated(433) xor estimated(434) xor estimated(435) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(28) <= estimated(112) xor estimated(113) xor estimated(114) xor estimated(115) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(29) <= estimated(368) xor estimated(369) xor estimated(370) xor estimated(371) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(30) <= estimated(240) xor estimated(241) xor estimated(242) xor estimated(243) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(31) <= estimated(496) xor estimated(497) xor estimated(498) xor estimated(499) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(32) <= estimated(8) xor estimated(9) xor estimated(10) xor estimated(11) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(33) <= estimated(264) xor estimated(265) xor estimated(266) xor estimated(267) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(34) <= estimated(136) xor estimated(137) xor estimated(138) xor estimated(139) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(35) <= estimated(392) xor estimated(393) xor estimated(394) xor estimated(395) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(36) <= estimated(72) xor estimated(73) xor estimated(74) xor estimated(75) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(37) <= estimated(328) xor estimated(329) xor estimated(330) xor estimated(331) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(38) <= estimated(200) xor estimated(201) xor estimated(202) xor estimated(203) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(39) <= estimated(456) xor estimated(457) xor estimated(458) xor estimated(459) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(40) <= estimated(40) xor estimated(41) xor estimated(42) xor estimated(43) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(41) <= estimated(296) xor estimated(297) xor estimated(298) xor estimated(299) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(42) <= estimated(168) xor estimated(169) xor estimated(170) xor estimated(171) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(43) <= estimated(424) xor estimated(425) xor estimated(426) xor estimated(427) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(44) <= estimated(104) xor estimated(105) xor estimated(106) xor estimated(107) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(45) <= estimated(360) xor estimated(361) xor estimated(362) xor estimated(363) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(46) <= estimated(232) xor estimated(233) xor estimated(234) xor estimated(235) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(47) <= estimated(488) xor estimated(489) xor estimated(490) xor estimated(491) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(48) <= estimated(24) xor estimated(25) xor estimated(26) xor estimated(27) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(49) <= estimated(280) xor estimated(281) xor estimated(282) xor estimated(283) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(50) <= estimated(152) xor estimated(153) xor estimated(154) xor estimated(155) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(51) <= estimated(408) xor estimated(409) xor estimated(410) xor estimated(411) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(52) <= estimated(88) xor estimated(89) xor estimated(90) xor estimated(91) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(53) <= estimated(344) xor estimated(345) xor estimated(346) xor estimated(347) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(54) <= estimated(216) xor estimated(217) xor estimated(218) xor estimated(219) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(55) <= estimated(472) xor estimated(473) xor estimated(474) xor estimated(475) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(56) <= estimated(56) xor estimated(57) xor estimated(58) xor estimated(59) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(57) <= estimated(312) xor estimated(313) xor estimated(314) xor estimated(315) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(58) <= estimated(184) xor estimated(185) xor estimated(186) xor estimated(187) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(59) <= estimated(440) xor estimated(441) xor estimated(442) xor estimated(443) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(60) <= estimated(120) xor estimated(121) xor estimated(122) xor estimated(123) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(61) <= estimated(376) xor estimated(377) xor estimated(378) xor estimated(379) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(62) <= estimated(248) xor estimated(249) xor estimated(250) xor estimated(251) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(63) <= estimated(504) xor estimated(505) xor estimated(506) xor estimated(507) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(64) <= estimated(4) xor estimated(5) xor estimated(6) xor estimated(7) xor estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(65) <= estimated(260) xor estimated(261) xor estimated(262) xor estimated(263) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(66) <= estimated(132) xor estimated(133) xor estimated(134) xor estimated(135) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(67) <= estimated(388) xor estimated(389) xor estimated(390) xor estimated(391) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(68) <= estimated(68) xor estimated(69) xor estimated(70) xor estimated(71) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(69) <= estimated(324) xor estimated(325) xor estimated(326) xor estimated(327) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(70) <= estimated(196) xor estimated(197) xor estimated(198) xor estimated(199) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(71) <= estimated(452) xor estimated(453) xor estimated(454) xor estimated(455) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(72) <= estimated(36) xor estimated(37) xor estimated(38) xor estimated(39) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(73) <= estimated(292) xor estimated(293) xor estimated(294) xor estimated(295) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(74) <= estimated(164) xor estimated(165) xor estimated(166) xor estimated(167) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(75) <= estimated(420) xor estimated(421) xor estimated(422) xor estimated(423) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(76) <= estimated(100) xor estimated(101) xor estimated(102) xor estimated(103) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(77) <= estimated(356) xor estimated(357) xor estimated(358) xor estimated(359) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(78) <= estimated(228) xor estimated(229) xor estimated(230) xor estimated(231) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(79) <= estimated(484) xor estimated(485) xor estimated(486) xor estimated(487) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(80) <= estimated(20) xor estimated(21) xor estimated(22) xor estimated(23) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(81) <= estimated(276) xor estimated(277) xor estimated(278) xor estimated(279) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(82) <= estimated(148) xor estimated(149) xor estimated(150) xor estimated(151) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(83) <= estimated(404) xor estimated(405) xor estimated(406) xor estimated(407) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(84) <= estimated(84) xor estimated(85) xor estimated(86) xor estimated(87) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(85) <= estimated(340) xor estimated(341) xor estimated(342) xor estimated(343) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(86) <= estimated(212) xor estimated(213) xor estimated(214) xor estimated(215) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(87) <= estimated(468) xor estimated(469) xor estimated(470) xor estimated(471) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(88) <= estimated(52) xor estimated(53) xor estimated(54) xor estimated(55) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(89) <= estimated(308) xor estimated(309) xor estimated(310) xor estimated(311) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(90) <= estimated(180) xor estimated(181) xor estimated(182) xor estimated(183) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(91) <= estimated(436) xor estimated(437) xor estimated(438) xor estimated(439) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(92) <= estimated(116) xor estimated(117) xor estimated(118) xor estimated(119) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(93) <= estimated(372) xor estimated(373) xor estimated(374) xor estimated(375) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(94) <= estimated(244) xor estimated(245) xor estimated(246) xor estimated(247) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(95) <= estimated(500) xor estimated(501) xor estimated(502) xor estimated(503) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(96) <= estimated(12) xor estimated(13) xor estimated(14) xor estimated(15) xor estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(97) <= estimated(268) xor estimated(269) xor estimated(270) xor estimated(271) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(98) <= estimated(140) xor estimated(141) xor estimated(142) xor estimated(143) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(99) <= estimated(396) xor estimated(397) xor estimated(398) xor estimated(399) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(100) <= estimated(76) xor estimated(77) xor estimated(78) xor estimated(79) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(101) <= estimated(332) xor estimated(333) xor estimated(334) xor estimated(335) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(102) <= estimated(204) xor estimated(205) xor estimated(206) xor estimated(207) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(103) <= estimated(460) xor estimated(461) xor estimated(462) xor estimated(463) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(104) <= estimated(44) xor estimated(45) xor estimated(46) xor estimated(47) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(105) <= estimated(300) xor estimated(301) xor estimated(302) xor estimated(303) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(106) <= estimated(172) xor estimated(173) xor estimated(174) xor estimated(175) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(107) <= estimated(428) xor estimated(429) xor estimated(430) xor estimated(431) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(108) <= estimated(108) xor estimated(109) xor estimated(110) xor estimated(111) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(109) <= estimated(364) xor estimated(365) xor estimated(366) xor estimated(367) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(110) <= estimated(236) xor estimated(237) xor estimated(238) xor estimated(239) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(111) <= estimated(492) xor estimated(493) xor estimated(494) xor estimated(495) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(112) <= estimated(28) xor estimated(29) xor estimated(30) xor estimated(31) xor estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(113) <= estimated(284) xor estimated(285) xor estimated(286) xor estimated(287) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(114) <= estimated(156) xor estimated(157) xor estimated(158) xor estimated(159) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(115) <= estimated(412) xor estimated(413) xor estimated(414) xor estimated(415) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(116) <= estimated(92) xor estimated(93) xor estimated(94) xor estimated(95) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(117) <= estimated(348) xor estimated(349) xor estimated(350) xor estimated(351) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(118) <= estimated(220) xor estimated(221) xor estimated(222) xor estimated(223) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(119) <= estimated(476) xor estimated(477) xor estimated(478) xor estimated(479) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(120) <= estimated(60) xor estimated(61) xor estimated(62) xor estimated(63) xor estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(121) <= estimated(316) xor estimated(317) xor estimated(318) xor estimated(319) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(122) <= estimated(188) xor estimated(189) xor estimated(190) xor estimated(191) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(123) <= estimated(444) xor estimated(445) xor estimated(446) xor estimated(447) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(124) <= estimated(124) xor estimated(125) xor estimated(126) xor estimated(127) xor estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(125) <= estimated(380) xor estimated(381) xor estimated(382) xor estimated(383) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(126) <= estimated(252) xor estimated(253) xor estimated(254) xor estimated(255) xor estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(127) <= estimated(508) xor estimated(509) xor estimated(510) xor estimated(511);
partial_sums(10)(128) <= estimated(2) xor estimated(3) xor estimated(6) xor estimated(7) xor estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(129) <= estimated(258) xor estimated(259) xor estimated(262) xor estimated(263) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(130) <= estimated(130) xor estimated(131) xor estimated(134) xor estimated(135) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(131) <= estimated(386) xor estimated(387) xor estimated(390) xor estimated(391) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(132) <= estimated(66) xor estimated(67) xor estimated(70) xor estimated(71) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(133) <= estimated(322) xor estimated(323) xor estimated(326) xor estimated(327) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(134) <= estimated(194) xor estimated(195) xor estimated(198) xor estimated(199) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(135) <= estimated(450) xor estimated(451) xor estimated(454) xor estimated(455) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(136) <= estimated(34) xor estimated(35) xor estimated(38) xor estimated(39) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(137) <= estimated(290) xor estimated(291) xor estimated(294) xor estimated(295) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(138) <= estimated(162) xor estimated(163) xor estimated(166) xor estimated(167) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(139) <= estimated(418) xor estimated(419) xor estimated(422) xor estimated(423) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(140) <= estimated(98) xor estimated(99) xor estimated(102) xor estimated(103) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(141) <= estimated(354) xor estimated(355) xor estimated(358) xor estimated(359) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(142) <= estimated(226) xor estimated(227) xor estimated(230) xor estimated(231) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(143) <= estimated(482) xor estimated(483) xor estimated(486) xor estimated(487) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(144) <= estimated(18) xor estimated(19) xor estimated(22) xor estimated(23) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(145) <= estimated(274) xor estimated(275) xor estimated(278) xor estimated(279) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(146) <= estimated(146) xor estimated(147) xor estimated(150) xor estimated(151) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(147) <= estimated(402) xor estimated(403) xor estimated(406) xor estimated(407) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(148) <= estimated(82) xor estimated(83) xor estimated(86) xor estimated(87) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(149) <= estimated(338) xor estimated(339) xor estimated(342) xor estimated(343) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(150) <= estimated(210) xor estimated(211) xor estimated(214) xor estimated(215) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(151) <= estimated(466) xor estimated(467) xor estimated(470) xor estimated(471) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(152) <= estimated(50) xor estimated(51) xor estimated(54) xor estimated(55) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(153) <= estimated(306) xor estimated(307) xor estimated(310) xor estimated(311) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(154) <= estimated(178) xor estimated(179) xor estimated(182) xor estimated(183) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(155) <= estimated(434) xor estimated(435) xor estimated(438) xor estimated(439) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(156) <= estimated(114) xor estimated(115) xor estimated(118) xor estimated(119) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(157) <= estimated(370) xor estimated(371) xor estimated(374) xor estimated(375) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(158) <= estimated(242) xor estimated(243) xor estimated(246) xor estimated(247) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(159) <= estimated(498) xor estimated(499) xor estimated(502) xor estimated(503) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(160) <= estimated(10) xor estimated(11) xor estimated(14) xor estimated(15) xor estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(161) <= estimated(266) xor estimated(267) xor estimated(270) xor estimated(271) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(162) <= estimated(138) xor estimated(139) xor estimated(142) xor estimated(143) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(163) <= estimated(394) xor estimated(395) xor estimated(398) xor estimated(399) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(164) <= estimated(74) xor estimated(75) xor estimated(78) xor estimated(79) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(165) <= estimated(330) xor estimated(331) xor estimated(334) xor estimated(335) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(166) <= estimated(202) xor estimated(203) xor estimated(206) xor estimated(207) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(167) <= estimated(458) xor estimated(459) xor estimated(462) xor estimated(463) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(168) <= estimated(42) xor estimated(43) xor estimated(46) xor estimated(47) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(169) <= estimated(298) xor estimated(299) xor estimated(302) xor estimated(303) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(170) <= estimated(170) xor estimated(171) xor estimated(174) xor estimated(175) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(171) <= estimated(426) xor estimated(427) xor estimated(430) xor estimated(431) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(172) <= estimated(106) xor estimated(107) xor estimated(110) xor estimated(111) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(173) <= estimated(362) xor estimated(363) xor estimated(366) xor estimated(367) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(174) <= estimated(234) xor estimated(235) xor estimated(238) xor estimated(239) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(175) <= estimated(490) xor estimated(491) xor estimated(494) xor estimated(495) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(176) <= estimated(26) xor estimated(27) xor estimated(30) xor estimated(31) xor estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(177) <= estimated(282) xor estimated(283) xor estimated(286) xor estimated(287) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(178) <= estimated(154) xor estimated(155) xor estimated(158) xor estimated(159) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(179) <= estimated(410) xor estimated(411) xor estimated(414) xor estimated(415) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(180) <= estimated(90) xor estimated(91) xor estimated(94) xor estimated(95) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(181) <= estimated(346) xor estimated(347) xor estimated(350) xor estimated(351) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(182) <= estimated(218) xor estimated(219) xor estimated(222) xor estimated(223) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(183) <= estimated(474) xor estimated(475) xor estimated(478) xor estimated(479) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(184) <= estimated(58) xor estimated(59) xor estimated(62) xor estimated(63) xor estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(185) <= estimated(314) xor estimated(315) xor estimated(318) xor estimated(319) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(186) <= estimated(186) xor estimated(187) xor estimated(190) xor estimated(191) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(187) <= estimated(442) xor estimated(443) xor estimated(446) xor estimated(447) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(188) <= estimated(122) xor estimated(123) xor estimated(126) xor estimated(127) xor estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(189) <= estimated(378) xor estimated(379) xor estimated(382) xor estimated(383) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(190) <= estimated(250) xor estimated(251) xor estimated(254) xor estimated(255) xor estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(191) <= estimated(506) xor estimated(507) xor estimated(510) xor estimated(511);
partial_sums(10)(192) <= estimated(6) xor estimated(7) xor estimated(14) xor estimated(15) xor estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(193) <= estimated(262) xor estimated(263) xor estimated(270) xor estimated(271) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(194) <= estimated(134) xor estimated(135) xor estimated(142) xor estimated(143) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(195) <= estimated(390) xor estimated(391) xor estimated(398) xor estimated(399) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(196) <= estimated(70) xor estimated(71) xor estimated(78) xor estimated(79) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(197) <= estimated(326) xor estimated(327) xor estimated(334) xor estimated(335) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(198) <= estimated(198) xor estimated(199) xor estimated(206) xor estimated(207) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(199) <= estimated(454) xor estimated(455) xor estimated(462) xor estimated(463) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(200) <= estimated(38) xor estimated(39) xor estimated(46) xor estimated(47) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(201) <= estimated(294) xor estimated(295) xor estimated(302) xor estimated(303) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(202) <= estimated(166) xor estimated(167) xor estimated(174) xor estimated(175) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(203) <= estimated(422) xor estimated(423) xor estimated(430) xor estimated(431) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(204) <= estimated(102) xor estimated(103) xor estimated(110) xor estimated(111) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(205) <= estimated(358) xor estimated(359) xor estimated(366) xor estimated(367) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(206) <= estimated(230) xor estimated(231) xor estimated(238) xor estimated(239) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(207) <= estimated(486) xor estimated(487) xor estimated(494) xor estimated(495) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(208) <= estimated(22) xor estimated(23) xor estimated(30) xor estimated(31) xor estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(209) <= estimated(278) xor estimated(279) xor estimated(286) xor estimated(287) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(210) <= estimated(150) xor estimated(151) xor estimated(158) xor estimated(159) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(211) <= estimated(406) xor estimated(407) xor estimated(414) xor estimated(415) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(212) <= estimated(86) xor estimated(87) xor estimated(94) xor estimated(95) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(213) <= estimated(342) xor estimated(343) xor estimated(350) xor estimated(351) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(214) <= estimated(214) xor estimated(215) xor estimated(222) xor estimated(223) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(215) <= estimated(470) xor estimated(471) xor estimated(478) xor estimated(479) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(216) <= estimated(54) xor estimated(55) xor estimated(62) xor estimated(63) xor estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(217) <= estimated(310) xor estimated(311) xor estimated(318) xor estimated(319) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(218) <= estimated(182) xor estimated(183) xor estimated(190) xor estimated(191) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(219) <= estimated(438) xor estimated(439) xor estimated(446) xor estimated(447) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(220) <= estimated(118) xor estimated(119) xor estimated(126) xor estimated(127) xor estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(221) <= estimated(374) xor estimated(375) xor estimated(382) xor estimated(383) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(222) <= estimated(246) xor estimated(247) xor estimated(254) xor estimated(255) xor estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(223) <= estimated(502) xor estimated(503) xor estimated(510) xor estimated(511);
partial_sums(10)(224) <= estimated(14) xor estimated(15) xor estimated(30) xor estimated(31) xor estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(270) xor estimated(271) xor estimated(286) xor estimated(287) xor estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(398) xor estimated(399) xor estimated(414) xor estimated(415) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(225) <= estimated(270) xor estimated(271) xor estimated(286) xor estimated(287) xor estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(398) xor estimated(399) xor estimated(414) xor estimated(415) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(226) <= estimated(142) xor estimated(143) xor estimated(158) xor estimated(159) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(398) xor estimated(399) xor estimated(414) xor estimated(415) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(227) <= estimated(398) xor estimated(399) xor estimated(414) xor estimated(415) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(228) <= estimated(78) xor estimated(79) xor estimated(94) xor estimated(95) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(229) <= estimated(334) xor estimated(335) xor estimated(350) xor estimated(351) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(230) <= estimated(206) xor estimated(207) xor estimated(222) xor estimated(223) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(231) <= estimated(462) xor estimated(463) xor estimated(478) xor estimated(479) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(232) <= estimated(46) xor estimated(47) xor estimated(62) xor estimated(63) xor estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(233) <= estimated(302) xor estimated(303) xor estimated(318) xor estimated(319) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(234) <= estimated(174) xor estimated(175) xor estimated(190) xor estimated(191) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(235) <= estimated(430) xor estimated(431) xor estimated(446) xor estimated(447) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(236) <= estimated(110) xor estimated(111) xor estimated(126) xor estimated(127) xor estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(237) <= estimated(366) xor estimated(367) xor estimated(382) xor estimated(383) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(238) <= estimated(238) xor estimated(239) xor estimated(254) xor estimated(255) xor estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(239) <= estimated(494) xor estimated(495) xor estimated(510) xor estimated(511);
partial_sums(10)(240) <= estimated(30) xor estimated(31) xor estimated(62) xor estimated(63) xor estimated(94) xor estimated(95) xor estimated(126) xor estimated(127) xor estimated(158) xor estimated(159) xor estimated(190) xor estimated(191) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255) xor estimated(286) xor estimated(287) xor estimated(318) xor estimated(319) xor estimated(350) xor estimated(351) xor estimated(382) xor estimated(383) xor estimated(414) xor estimated(415) xor estimated(446) xor estimated(447) xor estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(241) <= estimated(286) xor estimated(287) xor estimated(318) xor estimated(319) xor estimated(350) xor estimated(351) xor estimated(382) xor estimated(383) xor estimated(414) xor estimated(415) xor estimated(446) xor estimated(447) xor estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(242) <= estimated(158) xor estimated(159) xor estimated(190) xor estimated(191) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255) xor estimated(414) xor estimated(415) xor estimated(446) xor estimated(447) xor estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(243) <= estimated(414) xor estimated(415) xor estimated(446) xor estimated(447) xor estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(244) <= estimated(94) xor estimated(95) xor estimated(126) xor estimated(127) xor estimated(222) xor estimated(223) xor estimated(254) xor estimated(255) xor estimated(350) xor estimated(351) xor estimated(382) xor estimated(383) xor estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(245) <= estimated(350) xor estimated(351) xor estimated(382) xor estimated(383) xor estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(246) <= estimated(222) xor estimated(223) xor estimated(254) xor estimated(255) xor estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(247) <= estimated(478) xor estimated(479) xor estimated(510) xor estimated(511);
partial_sums(10)(248) <= estimated(62) xor estimated(63) xor estimated(126) xor estimated(127) xor estimated(190) xor estimated(191) xor estimated(254) xor estimated(255) xor estimated(318) xor estimated(319) xor estimated(382) xor estimated(383) xor estimated(446) xor estimated(447) xor estimated(510) xor estimated(511);
partial_sums(10)(249) <= estimated(318) xor estimated(319) xor estimated(382) xor estimated(383) xor estimated(446) xor estimated(447) xor estimated(510) xor estimated(511);
partial_sums(10)(250) <= estimated(190) xor estimated(191) xor estimated(254) xor estimated(255) xor estimated(446) xor estimated(447) xor estimated(510) xor estimated(511);
partial_sums(10)(251) <= estimated(446) xor estimated(447) xor estimated(510) xor estimated(511);
partial_sums(10)(252) <= estimated(126) xor estimated(127) xor estimated(254) xor estimated(255) xor estimated(382) xor estimated(383) xor estimated(510) xor estimated(511);
partial_sums(10)(253) <= estimated(382) xor estimated(383) xor estimated(510) xor estimated(511);
partial_sums(10)(254) <= estimated(254) xor estimated(255) xor estimated(510) xor estimated(511);
partial_sums(10)(255) <= estimated(510) xor estimated(511);
partial_sums(10)(256) <= estimated(1) xor estimated(3) xor estimated(5) xor estimated(7) xor estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(257) <= estimated(257) xor estimated(259) xor estimated(261) xor estimated(263) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(258) <= estimated(129) xor estimated(131) xor estimated(133) xor estimated(135) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(259) <= estimated(385) xor estimated(387) xor estimated(389) xor estimated(391) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(260) <= estimated(65) xor estimated(67) xor estimated(69) xor estimated(71) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(261) <= estimated(321) xor estimated(323) xor estimated(325) xor estimated(327) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(262) <= estimated(193) xor estimated(195) xor estimated(197) xor estimated(199) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(263) <= estimated(449) xor estimated(451) xor estimated(453) xor estimated(455) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(264) <= estimated(33) xor estimated(35) xor estimated(37) xor estimated(39) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(265) <= estimated(289) xor estimated(291) xor estimated(293) xor estimated(295) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(266) <= estimated(161) xor estimated(163) xor estimated(165) xor estimated(167) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(267) <= estimated(417) xor estimated(419) xor estimated(421) xor estimated(423) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(268) <= estimated(97) xor estimated(99) xor estimated(101) xor estimated(103) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(269) <= estimated(353) xor estimated(355) xor estimated(357) xor estimated(359) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(270) <= estimated(225) xor estimated(227) xor estimated(229) xor estimated(231) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(271) <= estimated(481) xor estimated(483) xor estimated(485) xor estimated(487) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(272) <= estimated(17) xor estimated(19) xor estimated(21) xor estimated(23) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(273) <= estimated(273) xor estimated(275) xor estimated(277) xor estimated(279) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(274) <= estimated(145) xor estimated(147) xor estimated(149) xor estimated(151) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(275) <= estimated(401) xor estimated(403) xor estimated(405) xor estimated(407) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(276) <= estimated(81) xor estimated(83) xor estimated(85) xor estimated(87) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(277) <= estimated(337) xor estimated(339) xor estimated(341) xor estimated(343) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(278) <= estimated(209) xor estimated(211) xor estimated(213) xor estimated(215) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(279) <= estimated(465) xor estimated(467) xor estimated(469) xor estimated(471) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(280) <= estimated(49) xor estimated(51) xor estimated(53) xor estimated(55) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(281) <= estimated(305) xor estimated(307) xor estimated(309) xor estimated(311) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(282) <= estimated(177) xor estimated(179) xor estimated(181) xor estimated(183) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(283) <= estimated(433) xor estimated(435) xor estimated(437) xor estimated(439) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(284) <= estimated(113) xor estimated(115) xor estimated(117) xor estimated(119) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(285) <= estimated(369) xor estimated(371) xor estimated(373) xor estimated(375) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(286) <= estimated(241) xor estimated(243) xor estimated(245) xor estimated(247) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(287) <= estimated(497) xor estimated(499) xor estimated(501) xor estimated(503) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(288) <= estimated(9) xor estimated(11) xor estimated(13) xor estimated(15) xor estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(289) <= estimated(265) xor estimated(267) xor estimated(269) xor estimated(271) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(290) <= estimated(137) xor estimated(139) xor estimated(141) xor estimated(143) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(291) <= estimated(393) xor estimated(395) xor estimated(397) xor estimated(399) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(292) <= estimated(73) xor estimated(75) xor estimated(77) xor estimated(79) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(293) <= estimated(329) xor estimated(331) xor estimated(333) xor estimated(335) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(294) <= estimated(201) xor estimated(203) xor estimated(205) xor estimated(207) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(295) <= estimated(457) xor estimated(459) xor estimated(461) xor estimated(463) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(296) <= estimated(41) xor estimated(43) xor estimated(45) xor estimated(47) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(297) <= estimated(297) xor estimated(299) xor estimated(301) xor estimated(303) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(298) <= estimated(169) xor estimated(171) xor estimated(173) xor estimated(175) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(299) <= estimated(425) xor estimated(427) xor estimated(429) xor estimated(431) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(300) <= estimated(105) xor estimated(107) xor estimated(109) xor estimated(111) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(301) <= estimated(361) xor estimated(363) xor estimated(365) xor estimated(367) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(302) <= estimated(233) xor estimated(235) xor estimated(237) xor estimated(239) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(303) <= estimated(489) xor estimated(491) xor estimated(493) xor estimated(495) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(304) <= estimated(25) xor estimated(27) xor estimated(29) xor estimated(31) xor estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(305) <= estimated(281) xor estimated(283) xor estimated(285) xor estimated(287) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(306) <= estimated(153) xor estimated(155) xor estimated(157) xor estimated(159) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(307) <= estimated(409) xor estimated(411) xor estimated(413) xor estimated(415) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(308) <= estimated(89) xor estimated(91) xor estimated(93) xor estimated(95) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(309) <= estimated(345) xor estimated(347) xor estimated(349) xor estimated(351) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(310) <= estimated(217) xor estimated(219) xor estimated(221) xor estimated(223) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(311) <= estimated(473) xor estimated(475) xor estimated(477) xor estimated(479) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(312) <= estimated(57) xor estimated(59) xor estimated(61) xor estimated(63) xor estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(313) <= estimated(313) xor estimated(315) xor estimated(317) xor estimated(319) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(314) <= estimated(185) xor estimated(187) xor estimated(189) xor estimated(191) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(315) <= estimated(441) xor estimated(443) xor estimated(445) xor estimated(447) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(316) <= estimated(121) xor estimated(123) xor estimated(125) xor estimated(127) xor estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(317) <= estimated(377) xor estimated(379) xor estimated(381) xor estimated(383) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(318) <= estimated(249) xor estimated(251) xor estimated(253) xor estimated(255) xor estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(319) <= estimated(505) xor estimated(507) xor estimated(509) xor estimated(511);
partial_sums(10)(320) <= estimated(5) xor estimated(7) xor estimated(13) xor estimated(15) xor estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(321) <= estimated(261) xor estimated(263) xor estimated(269) xor estimated(271) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(322) <= estimated(133) xor estimated(135) xor estimated(141) xor estimated(143) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(323) <= estimated(389) xor estimated(391) xor estimated(397) xor estimated(399) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(324) <= estimated(69) xor estimated(71) xor estimated(77) xor estimated(79) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(325) <= estimated(325) xor estimated(327) xor estimated(333) xor estimated(335) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(326) <= estimated(197) xor estimated(199) xor estimated(205) xor estimated(207) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(327) <= estimated(453) xor estimated(455) xor estimated(461) xor estimated(463) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(328) <= estimated(37) xor estimated(39) xor estimated(45) xor estimated(47) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(329) <= estimated(293) xor estimated(295) xor estimated(301) xor estimated(303) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(330) <= estimated(165) xor estimated(167) xor estimated(173) xor estimated(175) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(331) <= estimated(421) xor estimated(423) xor estimated(429) xor estimated(431) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(332) <= estimated(101) xor estimated(103) xor estimated(109) xor estimated(111) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(333) <= estimated(357) xor estimated(359) xor estimated(365) xor estimated(367) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(334) <= estimated(229) xor estimated(231) xor estimated(237) xor estimated(239) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(335) <= estimated(485) xor estimated(487) xor estimated(493) xor estimated(495) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(336) <= estimated(21) xor estimated(23) xor estimated(29) xor estimated(31) xor estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(337) <= estimated(277) xor estimated(279) xor estimated(285) xor estimated(287) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(338) <= estimated(149) xor estimated(151) xor estimated(157) xor estimated(159) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(339) <= estimated(405) xor estimated(407) xor estimated(413) xor estimated(415) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(340) <= estimated(85) xor estimated(87) xor estimated(93) xor estimated(95) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(341) <= estimated(341) xor estimated(343) xor estimated(349) xor estimated(351) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(342) <= estimated(213) xor estimated(215) xor estimated(221) xor estimated(223) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(343) <= estimated(469) xor estimated(471) xor estimated(477) xor estimated(479) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(344) <= estimated(53) xor estimated(55) xor estimated(61) xor estimated(63) xor estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(345) <= estimated(309) xor estimated(311) xor estimated(317) xor estimated(319) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(346) <= estimated(181) xor estimated(183) xor estimated(189) xor estimated(191) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(347) <= estimated(437) xor estimated(439) xor estimated(445) xor estimated(447) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(348) <= estimated(117) xor estimated(119) xor estimated(125) xor estimated(127) xor estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(349) <= estimated(373) xor estimated(375) xor estimated(381) xor estimated(383) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(350) <= estimated(245) xor estimated(247) xor estimated(253) xor estimated(255) xor estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(351) <= estimated(501) xor estimated(503) xor estimated(509) xor estimated(511);
partial_sums(10)(352) <= estimated(13) xor estimated(15) xor estimated(29) xor estimated(31) xor estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(269) xor estimated(271) xor estimated(285) xor estimated(287) xor estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(397) xor estimated(399) xor estimated(413) xor estimated(415) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(353) <= estimated(269) xor estimated(271) xor estimated(285) xor estimated(287) xor estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(397) xor estimated(399) xor estimated(413) xor estimated(415) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(354) <= estimated(141) xor estimated(143) xor estimated(157) xor estimated(159) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(397) xor estimated(399) xor estimated(413) xor estimated(415) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(355) <= estimated(397) xor estimated(399) xor estimated(413) xor estimated(415) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(356) <= estimated(77) xor estimated(79) xor estimated(93) xor estimated(95) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(357) <= estimated(333) xor estimated(335) xor estimated(349) xor estimated(351) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(358) <= estimated(205) xor estimated(207) xor estimated(221) xor estimated(223) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(359) <= estimated(461) xor estimated(463) xor estimated(477) xor estimated(479) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(360) <= estimated(45) xor estimated(47) xor estimated(61) xor estimated(63) xor estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(361) <= estimated(301) xor estimated(303) xor estimated(317) xor estimated(319) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(362) <= estimated(173) xor estimated(175) xor estimated(189) xor estimated(191) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(363) <= estimated(429) xor estimated(431) xor estimated(445) xor estimated(447) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(364) <= estimated(109) xor estimated(111) xor estimated(125) xor estimated(127) xor estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(365) <= estimated(365) xor estimated(367) xor estimated(381) xor estimated(383) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(366) <= estimated(237) xor estimated(239) xor estimated(253) xor estimated(255) xor estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(367) <= estimated(493) xor estimated(495) xor estimated(509) xor estimated(511);
partial_sums(10)(368) <= estimated(29) xor estimated(31) xor estimated(61) xor estimated(63) xor estimated(93) xor estimated(95) xor estimated(125) xor estimated(127) xor estimated(157) xor estimated(159) xor estimated(189) xor estimated(191) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255) xor estimated(285) xor estimated(287) xor estimated(317) xor estimated(319) xor estimated(349) xor estimated(351) xor estimated(381) xor estimated(383) xor estimated(413) xor estimated(415) xor estimated(445) xor estimated(447) xor estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(369) <= estimated(285) xor estimated(287) xor estimated(317) xor estimated(319) xor estimated(349) xor estimated(351) xor estimated(381) xor estimated(383) xor estimated(413) xor estimated(415) xor estimated(445) xor estimated(447) xor estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(370) <= estimated(157) xor estimated(159) xor estimated(189) xor estimated(191) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255) xor estimated(413) xor estimated(415) xor estimated(445) xor estimated(447) xor estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(371) <= estimated(413) xor estimated(415) xor estimated(445) xor estimated(447) xor estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(372) <= estimated(93) xor estimated(95) xor estimated(125) xor estimated(127) xor estimated(221) xor estimated(223) xor estimated(253) xor estimated(255) xor estimated(349) xor estimated(351) xor estimated(381) xor estimated(383) xor estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(373) <= estimated(349) xor estimated(351) xor estimated(381) xor estimated(383) xor estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(374) <= estimated(221) xor estimated(223) xor estimated(253) xor estimated(255) xor estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(375) <= estimated(477) xor estimated(479) xor estimated(509) xor estimated(511);
partial_sums(10)(376) <= estimated(61) xor estimated(63) xor estimated(125) xor estimated(127) xor estimated(189) xor estimated(191) xor estimated(253) xor estimated(255) xor estimated(317) xor estimated(319) xor estimated(381) xor estimated(383) xor estimated(445) xor estimated(447) xor estimated(509) xor estimated(511);
partial_sums(10)(377) <= estimated(317) xor estimated(319) xor estimated(381) xor estimated(383) xor estimated(445) xor estimated(447) xor estimated(509) xor estimated(511);
partial_sums(10)(378) <= estimated(189) xor estimated(191) xor estimated(253) xor estimated(255) xor estimated(445) xor estimated(447) xor estimated(509) xor estimated(511);
partial_sums(10)(379) <= estimated(445) xor estimated(447) xor estimated(509) xor estimated(511);
partial_sums(10)(380) <= estimated(125) xor estimated(127) xor estimated(253) xor estimated(255) xor estimated(381) xor estimated(383) xor estimated(509) xor estimated(511);
partial_sums(10)(381) <= estimated(381) xor estimated(383) xor estimated(509) xor estimated(511);
partial_sums(10)(382) <= estimated(253) xor estimated(255) xor estimated(509) xor estimated(511);
partial_sums(10)(383) <= estimated(509) xor estimated(511);
partial_sums(10)(384) <= estimated(3) xor estimated(7) xor estimated(11) xor estimated(15) xor estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(385) <= estimated(259) xor estimated(263) xor estimated(267) xor estimated(271) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(386) <= estimated(131) xor estimated(135) xor estimated(139) xor estimated(143) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(387) <= estimated(387) xor estimated(391) xor estimated(395) xor estimated(399) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(388) <= estimated(67) xor estimated(71) xor estimated(75) xor estimated(79) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(389) <= estimated(323) xor estimated(327) xor estimated(331) xor estimated(335) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(390) <= estimated(195) xor estimated(199) xor estimated(203) xor estimated(207) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(391) <= estimated(451) xor estimated(455) xor estimated(459) xor estimated(463) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(392) <= estimated(35) xor estimated(39) xor estimated(43) xor estimated(47) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(393) <= estimated(291) xor estimated(295) xor estimated(299) xor estimated(303) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(394) <= estimated(163) xor estimated(167) xor estimated(171) xor estimated(175) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(395) <= estimated(419) xor estimated(423) xor estimated(427) xor estimated(431) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(396) <= estimated(99) xor estimated(103) xor estimated(107) xor estimated(111) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(397) <= estimated(355) xor estimated(359) xor estimated(363) xor estimated(367) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(398) <= estimated(227) xor estimated(231) xor estimated(235) xor estimated(239) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(399) <= estimated(483) xor estimated(487) xor estimated(491) xor estimated(495) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(400) <= estimated(19) xor estimated(23) xor estimated(27) xor estimated(31) xor estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(401) <= estimated(275) xor estimated(279) xor estimated(283) xor estimated(287) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(402) <= estimated(147) xor estimated(151) xor estimated(155) xor estimated(159) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(403) <= estimated(403) xor estimated(407) xor estimated(411) xor estimated(415) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(404) <= estimated(83) xor estimated(87) xor estimated(91) xor estimated(95) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(405) <= estimated(339) xor estimated(343) xor estimated(347) xor estimated(351) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(406) <= estimated(211) xor estimated(215) xor estimated(219) xor estimated(223) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(407) <= estimated(467) xor estimated(471) xor estimated(475) xor estimated(479) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(408) <= estimated(51) xor estimated(55) xor estimated(59) xor estimated(63) xor estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(409) <= estimated(307) xor estimated(311) xor estimated(315) xor estimated(319) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(410) <= estimated(179) xor estimated(183) xor estimated(187) xor estimated(191) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(411) <= estimated(435) xor estimated(439) xor estimated(443) xor estimated(447) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(412) <= estimated(115) xor estimated(119) xor estimated(123) xor estimated(127) xor estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(413) <= estimated(371) xor estimated(375) xor estimated(379) xor estimated(383) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(414) <= estimated(243) xor estimated(247) xor estimated(251) xor estimated(255) xor estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(415) <= estimated(499) xor estimated(503) xor estimated(507) xor estimated(511);
partial_sums(10)(416) <= estimated(11) xor estimated(15) xor estimated(27) xor estimated(31) xor estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(267) xor estimated(271) xor estimated(283) xor estimated(287) xor estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(395) xor estimated(399) xor estimated(411) xor estimated(415) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(417) <= estimated(267) xor estimated(271) xor estimated(283) xor estimated(287) xor estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(395) xor estimated(399) xor estimated(411) xor estimated(415) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(418) <= estimated(139) xor estimated(143) xor estimated(155) xor estimated(159) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(395) xor estimated(399) xor estimated(411) xor estimated(415) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(419) <= estimated(395) xor estimated(399) xor estimated(411) xor estimated(415) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(420) <= estimated(75) xor estimated(79) xor estimated(91) xor estimated(95) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(421) <= estimated(331) xor estimated(335) xor estimated(347) xor estimated(351) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(422) <= estimated(203) xor estimated(207) xor estimated(219) xor estimated(223) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(423) <= estimated(459) xor estimated(463) xor estimated(475) xor estimated(479) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(424) <= estimated(43) xor estimated(47) xor estimated(59) xor estimated(63) xor estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(425) <= estimated(299) xor estimated(303) xor estimated(315) xor estimated(319) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(426) <= estimated(171) xor estimated(175) xor estimated(187) xor estimated(191) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(427) <= estimated(427) xor estimated(431) xor estimated(443) xor estimated(447) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(428) <= estimated(107) xor estimated(111) xor estimated(123) xor estimated(127) xor estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(429) <= estimated(363) xor estimated(367) xor estimated(379) xor estimated(383) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(430) <= estimated(235) xor estimated(239) xor estimated(251) xor estimated(255) xor estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(431) <= estimated(491) xor estimated(495) xor estimated(507) xor estimated(511);
partial_sums(10)(432) <= estimated(27) xor estimated(31) xor estimated(59) xor estimated(63) xor estimated(91) xor estimated(95) xor estimated(123) xor estimated(127) xor estimated(155) xor estimated(159) xor estimated(187) xor estimated(191) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255) xor estimated(283) xor estimated(287) xor estimated(315) xor estimated(319) xor estimated(347) xor estimated(351) xor estimated(379) xor estimated(383) xor estimated(411) xor estimated(415) xor estimated(443) xor estimated(447) xor estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(433) <= estimated(283) xor estimated(287) xor estimated(315) xor estimated(319) xor estimated(347) xor estimated(351) xor estimated(379) xor estimated(383) xor estimated(411) xor estimated(415) xor estimated(443) xor estimated(447) xor estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(434) <= estimated(155) xor estimated(159) xor estimated(187) xor estimated(191) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255) xor estimated(411) xor estimated(415) xor estimated(443) xor estimated(447) xor estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(435) <= estimated(411) xor estimated(415) xor estimated(443) xor estimated(447) xor estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(436) <= estimated(91) xor estimated(95) xor estimated(123) xor estimated(127) xor estimated(219) xor estimated(223) xor estimated(251) xor estimated(255) xor estimated(347) xor estimated(351) xor estimated(379) xor estimated(383) xor estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(437) <= estimated(347) xor estimated(351) xor estimated(379) xor estimated(383) xor estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(438) <= estimated(219) xor estimated(223) xor estimated(251) xor estimated(255) xor estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(439) <= estimated(475) xor estimated(479) xor estimated(507) xor estimated(511);
partial_sums(10)(440) <= estimated(59) xor estimated(63) xor estimated(123) xor estimated(127) xor estimated(187) xor estimated(191) xor estimated(251) xor estimated(255) xor estimated(315) xor estimated(319) xor estimated(379) xor estimated(383) xor estimated(443) xor estimated(447) xor estimated(507) xor estimated(511);
partial_sums(10)(441) <= estimated(315) xor estimated(319) xor estimated(379) xor estimated(383) xor estimated(443) xor estimated(447) xor estimated(507) xor estimated(511);
partial_sums(10)(442) <= estimated(187) xor estimated(191) xor estimated(251) xor estimated(255) xor estimated(443) xor estimated(447) xor estimated(507) xor estimated(511);
partial_sums(10)(443) <= estimated(443) xor estimated(447) xor estimated(507) xor estimated(511);
partial_sums(10)(444) <= estimated(123) xor estimated(127) xor estimated(251) xor estimated(255) xor estimated(379) xor estimated(383) xor estimated(507) xor estimated(511);
partial_sums(10)(445) <= estimated(379) xor estimated(383) xor estimated(507) xor estimated(511);
partial_sums(10)(446) <= estimated(251) xor estimated(255) xor estimated(507) xor estimated(511);
partial_sums(10)(447) <= estimated(507) xor estimated(511);
partial_sums(10)(448) <= estimated(7) xor estimated(15) xor estimated(23) xor estimated(31) xor estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(263) xor estimated(271) xor estimated(279) xor estimated(287) xor estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(391) xor estimated(399) xor estimated(407) xor estimated(415) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(449) <= estimated(263) xor estimated(271) xor estimated(279) xor estimated(287) xor estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(391) xor estimated(399) xor estimated(407) xor estimated(415) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(450) <= estimated(135) xor estimated(143) xor estimated(151) xor estimated(159) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(391) xor estimated(399) xor estimated(407) xor estimated(415) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(451) <= estimated(391) xor estimated(399) xor estimated(407) xor estimated(415) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(452) <= estimated(71) xor estimated(79) xor estimated(87) xor estimated(95) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(453) <= estimated(327) xor estimated(335) xor estimated(343) xor estimated(351) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(454) <= estimated(199) xor estimated(207) xor estimated(215) xor estimated(223) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(455) <= estimated(455) xor estimated(463) xor estimated(471) xor estimated(479) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(456) <= estimated(39) xor estimated(47) xor estimated(55) xor estimated(63) xor estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(457) <= estimated(295) xor estimated(303) xor estimated(311) xor estimated(319) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(458) <= estimated(167) xor estimated(175) xor estimated(183) xor estimated(191) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(459) <= estimated(423) xor estimated(431) xor estimated(439) xor estimated(447) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(460) <= estimated(103) xor estimated(111) xor estimated(119) xor estimated(127) xor estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(461) <= estimated(359) xor estimated(367) xor estimated(375) xor estimated(383) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(462) <= estimated(231) xor estimated(239) xor estimated(247) xor estimated(255) xor estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(463) <= estimated(487) xor estimated(495) xor estimated(503) xor estimated(511);
partial_sums(10)(464) <= estimated(23) xor estimated(31) xor estimated(55) xor estimated(63) xor estimated(87) xor estimated(95) xor estimated(119) xor estimated(127) xor estimated(151) xor estimated(159) xor estimated(183) xor estimated(191) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255) xor estimated(279) xor estimated(287) xor estimated(311) xor estimated(319) xor estimated(343) xor estimated(351) xor estimated(375) xor estimated(383) xor estimated(407) xor estimated(415) xor estimated(439) xor estimated(447) xor estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(465) <= estimated(279) xor estimated(287) xor estimated(311) xor estimated(319) xor estimated(343) xor estimated(351) xor estimated(375) xor estimated(383) xor estimated(407) xor estimated(415) xor estimated(439) xor estimated(447) xor estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(466) <= estimated(151) xor estimated(159) xor estimated(183) xor estimated(191) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255) xor estimated(407) xor estimated(415) xor estimated(439) xor estimated(447) xor estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(467) <= estimated(407) xor estimated(415) xor estimated(439) xor estimated(447) xor estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(468) <= estimated(87) xor estimated(95) xor estimated(119) xor estimated(127) xor estimated(215) xor estimated(223) xor estimated(247) xor estimated(255) xor estimated(343) xor estimated(351) xor estimated(375) xor estimated(383) xor estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(469) <= estimated(343) xor estimated(351) xor estimated(375) xor estimated(383) xor estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(470) <= estimated(215) xor estimated(223) xor estimated(247) xor estimated(255) xor estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(471) <= estimated(471) xor estimated(479) xor estimated(503) xor estimated(511);
partial_sums(10)(472) <= estimated(55) xor estimated(63) xor estimated(119) xor estimated(127) xor estimated(183) xor estimated(191) xor estimated(247) xor estimated(255) xor estimated(311) xor estimated(319) xor estimated(375) xor estimated(383) xor estimated(439) xor estimated(447) xor estimated(503) xor estimated(511);
partial_sums(10)(473) <= estimated(311) xor estimated(319) xor estimated(375) xor estimated(383) xor estimated(439) xor estimated(447) xor estimated(503) xor estimated(511);
partial_sums(10)(474) <= estimated(183) xor estimated(191) xor estimated(247) xor estimated(255) xor estimated(439) xor estimated(447) xor estimated(503) xor estimated(511);
partial_sums(10)(475) <= estimated(439) xor estimated(447) xor estimated(503) xor estimated(511);
partial_sums(10)(476) <= estimated(119) xor estimated(127) xor estimated(247) xor estimated(255) xor estimated(375) xor estimated(383) xor estimated(503) xor estimated(511);
partial_sums(10)(477) <= estimated(375) xor estimated(383) xor estimated(503) xor estimated(511);
partial_sums(10)(478) <= estimated(247) xor estimated(255) xor estimated(503) xor estimated(511);
partial_sums(10)(479) <= estimated(503) xor estimated(511);
partial_sums(10)(480) <= estimated(15) xor estimated(31) xor estimated(47) xor estimated(63) xor estimated(79) xor estimated(95) xor estimated(111) xor estimated(127) xor estimated(143) xor estimated(159) xor estimated(175) xor estimated(191) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255) xor estimated(271) xor estimated(287) xor estimated(303) xor estimated(319) xor estimated(335) xor estimated(351) xor estimated(367) xor estimated(383) xor estimated(399) xor estimated(415) xor estimated(431) xor estimated(447) xor estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(481) <= estimated(271) xor estimated(287) xor estimated(303) xor estimated(319) xor estimated(335) xor estimated(351) xor estimated(367) xor estimated(383) xor estimated(399) xor estimated(415) xor estimated(431) xor estimated(447) xor estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(482) <= estimated(143) xor estimated(159) xor estimated(175) xor estimated(191) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255) xor estimated(399) xor estimated(415) xor estimated(431) xor estimated(447) xor estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(483) <= estimated(399) xor estimated(415) xor estimated(431) xor estimated(447) xor estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(484) <= estimated(79) xor estimated(95) xor estimated(111) xor estimated(127) xor estimated(207) xor estimated(223) xor estimated(239) xor estimated(255) xor estimated(335) xor estimated(351) xor estimated(367) xor estimated(383) xor estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(485) <= estimated(335) xor estimated(351) xor estimated(367) xor estimated(383) xor estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(486) <= estimated(207) xor estimated(223) xor estimated(239) xor estimated(255) xor estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(487) <= estimated(463) xor estimated(479) xor estimated(495) xor estimated(511);
partial_sums(10)(488) <= estimated(47) xor estimated(63) xor estimated(111) xor estimated(127) xor estimated(175) xor estimated(191) xor estimated(239) xor estimated(255) xor estimated(303) xor estimated(319) xor estimated(367) xor estimated(383) xor estimated(431) xor estimated(447) xor estimated(495) xor estimated(511);
partial_sums(10)(489) <= estimated(303) xor estimated(319) xor estimated(367) xor estimated(383) xor estimated(431) xor estimated(447) xor estimated(495) xor estimated(511);
partial_sums(10)(490) <= estimated(175) xor estimated(191) xor estimated(239) xor estimated(255) xor estimated(431) xor estimated(447) xor estimated(495) xor estimated(511);
partial_sums(10)(491) <= estimated(431) xor estimated(447) xor estimated(495) xor estimated(511);
partial_sums(10)(492) <= estimated(111) xor estimated(127) xor estimated(239) xor estimated(255) xor estimated(367) xor estimated(383) xor estimated(495) xor estimated(511);
partial_sums(10)(493) <= estimated(367) xor estimated(383) xor estimated(495) xor estimated(511);
partial_sums(10)(494) <= estimated(239) xor estimated(255) xor estimated(495) xor estimated(511);
partial_sums(10)(495) <= estimated(495) xor estimated(511);
partial_sums(10)(496) <= estimated(31) xor estimated(63) xor estimated(95) xor estimated(127) xor estimated(159) xor estimated(191) xor estimated(223) xor estimated(255) xor estimated(287) xor estimated(319) xor estimated(351) xor estimated(383) xor estimated(415) xor estimated(447) xor estimated(479) xor estimated(511);
partial_sums(10)(497) <= estimated(287) xor estimated(319) xor estimated(351) xor estimated(383) xor estimated(415) xor estimated(447) xor estimated(479) xor estimated(511);
partial_sums(10)(498) <= estimated(159) xor estimated(191) xor estimated(223) xor estimated(255) xor estimated(415) xor estimated(447) xor estimated(479) xor estimated(511);
partial_sums(10)(499) <= estimated(415) xor estimated(447) xor estimated(479) xor estimated(511);
partial_sums(10)(500) <= estimated(95) xor estimated(127) xor estimated(223) xor estimated(255) xor estimated(351) xor estimated(383) xor estimated(479) xor estimated(511);
partial_sums(10)(501) <= estimated(351) xor estimated(383) xor estimated(479) xor estimated(511);
partial_sums(10)(502) <= estimated(223) xor estimated(255) xor estimated(479) xor estimated(511);
partial_sums(10)(503) <= estimated(479) xor estimated(511);
partial_sums(10)(504) <= estimated(63) xor estimated(127) xor estimated(191) xor estimated(255) xor estimated(319) xor estimated(383) xor estimated(447) xor estimated(511);
partial_sums(10)(505) <= estimated(319) xor estimated(383) xor estimated(447) xor estimated(511);
partial_sums(10)(506) <= estimated(191) xor estimated(255) xor estimated(447) xor estimated(511);
partial_sums(10)(507) <= estimated(447) xor estimated(511);
partial_sums(10)(508) <= estimated(127) xor estimated(255) xor estimated(383) xor estimated(511);
partial_sums(10)(509) <= estimated(383) xor estimated(511);
partial_sums(10)(510) <= estimated(255) xor estimated(511);
partial_sums(10)(511) <= estimated(511);

end Behavioral;


----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:50:12 04/01/2016 
-- Design Name: 
-- Module Name:    Decoder512 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.all;
use work.MyPackage.all;
use IEEE.math_real.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Decoder512 is
    Port ( clk : in  STD_LOGIC;
           rst : in STD_LOGIC;
			  ce_inputs: in STD_LOGIC;
			  inputs : in data;
           outputs : out  STD_LOGIC_VECTOR (N/2-1 downto 0));
end Decoder512;

architecture Behavioral of Decoder512 is
	signal P: llr_2d := (others=>(others=>(others=> '0')));
	signal u : std_logic_vector(0 to N-2) := (others => '0');
	signal s: s_2d := (others=>(others=> '0'));
	signal ce_outputs : std_logic := '1';
begin

--Input Registers
GEN_REG_INPUT:
	for I in 0 to N-1 generate
		D_FF_gen: entity D_FF_gen generic map(width => fractional_part+integer_part)
											port map(clk => clk,
											rst => rst,
											ce => ce_inputs,
											d => inputs(I),
											q => P(stages)(I));
	end generate GEN_REG_INPUT;

-- STAGE 9
F90: entity F port map(lamdaA => P(9)(0),lamdaB => P(9)(1),lamdaOut => P(8)(0));
G91: entity G port map(lamdaA => P(9)(0),lamdaB => P(9)(1),s => s(9)(0),lamdaOut => P(8)(1));
F92: entity F port map(lamdaA => P(9)(2),lamdaB => P(9)(3),lamdaOut => P(8)(2));
G93: entity G port map(lamdaA => P(9)(2),lamdaB => P(9)(3),s => s(9)(1),lamdaOut => P(8)(3));
F94: entity F port map(lamdaA => P(9)(4),lamdaB => P(9)(5),lamdaOut => P(8)(4));
G95: entity G port map(lamdaA => P(9)(4),lamdaB => P(9)(5),s => s(9)(2),lamdaOut => P(8)(5));
F96: entity F port map(lamdaA => P(9)(6),lamdaB => P(9)(7),lamdaOut => P(8)(6));
G97: entity G port map(lamdaA => P(9)(6),lamdaB => P(9)(7),s => s(9)(3),lamdaOut => P(8)(7));
F98: entity F port map(lamdaA => P(9)(8),lamdaB => P(9)(9),lamdaOut => P(8)(8));
G99: entity G port map(lamdaA => P(9)(8),lamdaB => P(9)(9),s => s(9)(4),lamdaOut => P(8)(9));
F910: entity F port map(lamdaA => P(9)(10),lamdaB => P(9)(11),lamdaOut => P(8)(10));
G911: entity G port map(lamdaA => P(9)(10),lamdaB => P(9)(11),s => s(9)(5),lamdaOut => P(8)(11));
F912: entity F port map(lamdaA => P(9)(12),lamdaB => P(9)(13),lamdaOut => P(8)(12));
G913: entity G port map(lamdaA => P(9)(12),lamdaB => P(9)(13),s => s(9)(6),lamdaOut => P(8)(13));
F914: entity F port map(lamdaA => P(9)(14),lamdaB => P(9)(15),lamdaOut => P(8)(14));
G915: entity G port map(lamdaA => P(9)(14),lamdaB => P(9)(15),s => s(9)(7),lamdaOut => P(8)(15));
F916: entity F port map(lamdaA => P(9)(16),lamdaB => P(9)(17),lamdaOut => P(8)(16));
G917: entity G port map(lamdaA => P(9)(16),lamdaB => P(9)(17),s => s(9)(8),lamdaOut => P(8)(17));
F918: entity F port map(lamdaA => P(9)(18),lamdaB => P(9)(19),lamdaOut => P(8)(18));
G919: entity G port map(lamdaA => P(9)(18),lamdaB => P(9)(19),s => s(9)(9),lamdaOut => P(8)(19));
F920: entity F port map(lamdaA => P(9)(20),lamdaB => P(9)(21),lamdaOut => P(8)(20));
G921: entity G port map(lamdaA => P(9)(20),lamdaB => P(9)(21),s => s(9)(10),lamdaOut => P(8)(21));
F922: entity F port map(lamdaA => P(9)(22),lamdaB => P(9)(23),lamdaOut => P(8)(22));
G923: entity G port map(lamdaA => P(9)(22),lamdaB => P(9)(23),s => s(9)(11),lamdaOut => P(8)(23));
F924: entity F port map(lamdaA => P(9)(24),lamdaB => P(9)(25),lamdaOut => P(8)(24));
G925: entity G port map(lamdaA => P(9)(24),lamdaB => P(9)(25),s => s(9)(12),lamdaOut => P(8)(25));
F926: entity F port map(lamdaA => P(9)(26),lamdaB => P(9)(27),lamdaOut => P(8)(26));
G927: entity G port map(lamdaA => P(9)(26),lamdaB => P(9)(27),s => s(9)(13),lamdaOut => P(8)(27));
F928: entity F port map(lamdaA => P(9)(28),lamdaB => P(9)(29),lamdaOut => P(8)(28));
G929: entity G port map(lamdaA => P(9)(28),lamdaB => P(9)(29),s => s(9)(14),lamdaOut => P(8)(29));
F930: entity F port map(lamdaA => P(9)(30),lamdaB => P(9)(31),lamdaOut => P(8)(30));
G931: entity G port map(lamdaA => P(9)(30),lamdaB => P(9)(31),s => s(9)(15),lamdaOut => P(8)(31));
F932: entity F port map(lamdaA => P(9)(32),lamdaB => P(9)(33),lamdaOut => P(8)(32));
G933: entity G port map(lamdaA => P(9)(32),lamdaB => P(9)(33),s => s(9)(16),lamdaOut => P(8)(33));
F934: entity F port map(lamdaA => P(9)(34),lamdaB => P(9)(35),lamdaOut => P(8)(34));
G935: entity G port map(lamdaA => P(9)(34),lamdaB => P(9)(35),s => s(9)(17),lamdaOut => P(8)(35));
F936: entity F port map(lamdaA => P(9)(36),lamdaB => P(9)(37),lamdaOut => P(8)(36));
G937: entity G port map(lamdaA => P(9)(36),lamdaB => P(9)(37),s => s(9)(18),lamdaOut => P(8)(37));
F938: entity F port map(lamdaA => P(9)(38),lamdaB => P(9)(39),lamdaOut => P(8)(38));
G939: entity G port map(lamdaA => P(9)(38),lamdaB => P(9)(39),s => s(9)(19),lamdaOut => P(8)(39));
F940: entity F port map(lamdaA => P(9)(40),lamdaB => P(9)(41),lamdaOut => P(8)(40));
G941: entity G port map(lamdaA => P(9)(40),lamdaB => P(9)(41),s => s(9)(20),lamdaOut => P(8)(41));
F942: entity F port map(lamdaA => P(9)(42),lamdaB => P(9)(43),lamdaOut => P(8)(42));
G943: entity G port map(lamdaA => P(9)(42),lamdaB => P(9)(43),s => s(9)(21),lamdaOut => P(8)(43));
F944: entity F port map(lamdaA => P(9)(44),lamdaB => P(9)(45),lamdaOut => P(8)(44));
G945: entity G port map(lamdaA => P(9)(44),lamdaB => P(9)(45),s => s(9)(22),lamdaOut => P(8)(45));
F946: entity F port map(lamdaA => P(9)(46),lamdaB => P(9)(47),lamdaOut => P(8)(46));
G947: entity G port map(lamdaA => P(9)(46),lamdaB => P(9)(47),s => s(9)(23),lamdaOut => P(8)(47));
F948: entity F port map(lamdaA => P(9)(48),lamdaB => P(9)(49),lamdaOut => P(8)(48));
G949: entity G port map(lamdaA => P(9)(48),lamdaB => P(9)(49),s => s(9)(24),lamdaOut => P(8)(49));
F950: entity F port map(lamdaA => P(9)(50),lamdaB => P(9)(51),lamdaOut => P(8)(50));
G951: entity G port map(lamdaA => P(9)(50),lamdaB => P(9)(51),s => s(9)(25),lamdaOut => P(8)(51));
F952: entity F port map(lamdaA => P(9)(52),lamdaB => P(9)(53),lamdaOut => P(8)(52));
G953: entity G port map(lamdaA => P(9)(52),lamdaB => P(9)(53),s => s(9)(26),lamdaOut => P(8)(53));
F954: entity F port map(lamdaA => P(9)(54),lamdaB => P(9)(55),lamdaOut => P(8)(54));
G955: entity G port map(lamdaA => P(9)(54),lamdaB => P(9)(55),s => s(9)(27),lamdaOut => P(8)(55));
F956: entity F port map(lamdaA => P(9)(56),lamdaB => P(9)(57),lamdaOut => P(8)(56));
G957: entity G port map(lamdaA => P(9)(56),lamdaB => P(9)(57),s => s(9)(28),lamdaOut => P(8)(57));
F958: entity F port map(lamdaA => P(9)(58),lamdaB => P(9)(59),lamdaOut => P(8)(58));
G959: entity G port map(lamdaA => P(9)(58),lamdaB => P(9)(59),s => s(9)(29),lamdaOut => P(8)(59));
F960: entity F port map(lamdaA => P(9)(60),lamdaB => P(9)(61),lamdaOut => P(8)(60));
G961: entity G port map(lamdaA => P(9)(60),lamdaB => P(9)(61),s => s(9)(30),lamdaOut => P(8)(61));
F962: entity F port map(lamdaA => P(9)(62),lamdaB => P(9)(63),lamdaOut => P(8)(62));
G963: entity G port map(lamdaA => P(9)(62),lamdaB => P(9)(63),s => s(9)(31),lamdaOut => P(8)(63));
F964: entity F port map(lamdaA => P(9)(64),lamdaB => P(9)(65),lamdaOut => P(8)(64));
G965: entity G port map(lamdaA => P(9)(64),lamdaB => P(9)(65),s => s(9)(32),lamdaOut => P(8)(65));
F966: entity F port map(lamdaA => P(9)(66),lamdaB => P(9)(67),lamdaOut => P(8)(66));
G967: entity G port map(lamdaA => P(9)(66),lamdaB => P(9)(67),s => s(9)(33),lamdaOut => P(8)(67));
F968: entity F port map(lamdaA => P(9)(68),lamdaB => P(9)(69),lamdaOut => P(8)(68));
G969: entity G port map(lamdaA => P(9)(68),lamdaB => P(9)(69),s => s(9)(34),lamdaOut => P(8)(69));
F970: entity F port map(lamdaA => P(9)(70),lamdaB => P(9)(71),lamdaOut => P(8)(70));
G971: entity G port map(lamdaA => P(9)(70),lamdaB => P(9)(71),s => s(9)(35),lamdaOut => P(8)(71));
F972: entity F port map(lamdaA => P(9)(72),lamdaB => P(9)(73),lamdaOut => P(8)(72));
G973: entity G port map(lamdaA => P(9)(72),lamdaB => P(9)(73),s => s(9)(36),lamdaOut => P(8)(73));
F974: entity F port map(lamdaA => P(9)(74),lamdaB => P(9)(75),lamdaOut => P(8)(74));
G975: entity G port map(lamdaA => P(9)(74),lamdaB => P(9)(75),s => s(9)(37),lamdaOut => P(8)(75));
F976: entity F port map(lamdaA => P(9)(76),lamdaB => P(9)(77),lamdaOut => P(8)(76));
G977: entity G port map(lamdaA => P(9)(76),lamdaB => P(9)(77),s => s(9)(38),lamdaOut => P(8)(77));
F978: entity F port map(lamdaA => P(9)(78),lamdaB => P(9)(79),lamdaOut => P(8)(78));
G979: entity G port map(lamdaA => P(9)(78),lamdaB => P(9)(79),s => s(9)(39),lamdaOut => P(8)(79));
F980: entity F port map(lamdaA => P(9)(80),lamdaB => P(9)(81),lamdaOut => P(8)(80));
G981: entity G port map(lamdaA => P(9)(80),lamdaB => P(9)(81),s => s(9)(40),lamdaOut => P(8)(81));
F982: entity F port map(lamdaA => P(9)(82),lamdaB => P(9)(83),lamdaOut => P(8)(82));
G983: entity G port map(lamdaA => P(9)(82),lamdaB => P(9)(83),s => s(9)(41),lamdaOut => P(8)(83));
F984: entity F port map(lamdaA => P(9)(84),lamdaB => P(9)(85),lamdaOut => P(8)(84));
G985: entity G port map(lamdaA => P(9)(84),lamdaB => P(9)(85),s => s(9)(42),lamdaOut => P(8)(85));
F986: entity F port map(lamdaA => P(9)(86),lamdaB => P(9)(87),lamdaOut => P(8)(86));
G987: entity G port map(lamdaA => P(9)(86),lamdaB => P(9)(87),s => s(9)(43),lamdaOut => P(8)(87));
F988: entity F port map(lamdaA => P(9)(88),lamdaB => P(9)(89),lamdaOut => P(8)(88));
G989: entity G port map(lamdaA => P(9)(88),lamdaB => P(9)(89),s => s(9)(44),lamdaOut => P(8)(89));
F990: entity F port map(lamdaA => P(9)(90),lamdaB => P(9)(91),lamdaOut => P(8)(90));
G991: entity G port map(lamdaA => P(9)(90),lamdaB => P(9)(91),s => s(9)(45),lamdaOut => P(8)(91));
F992: entity F port map(lamdaA => P(9)(92),lamdaB => P(9)(93),lamdaOut => P(8)(92));
G993: entity G port map(lamdaA => P(9)(92),lamdaB => P(9)(93),s => s(9)(46),lamdaOut => P(8)(93));
F994: entity F port map(lamdaA => P(9)(94),lamdaB => P(9)(95),lamdaOut => P(8)(94));
G995: entity G port map(lamdaA => P(9)(94),lamdaB => P(9)(95),s => s(9)(47),lamdaOut => P(8)(95));
F996: entity F port map(lamdaA => P(9)(96),lamdaB => P(9)(97),lamdaOut => P(8)(96));
G997: entity G port map(lamdaA => P(9)(96),lamdaB => P(9)(97),s => s(9)(48),lamdaOut => P(8)(97));
F998: entity F port map(lamdaA => P(9)(98),lamdaB => P(9)(99),lamdaOut => P(8)(98));
G999: entity G port map(lamdaA => P(9)(98),lamdaB => P(9)(99),s => s(9)(49),lamdaOut => P(8)(99));
F9100: entity F port map(lamdaA => P(9)(100),lamdaB => P(9)(101),lamdaOut => P(8)(100));
G9101: entity G port map(lamdaA => P(9)(100),lamdaB => P(9)(101),s => s(9)(50),lamdaOut => P(8)(101));
F9102: entity F port map(lamdaA => P(9)(102),lamdaB => P(9)(103),lamdaOut => P(8)(102));
G9103: entity G port map(lamdaA => P(9)(102),lamdaB => P(9)(103),s => s(9)(51),lamdaOut => P(8)(103));
F9104: entity F port map(lamdaA => P(9)(104),lamdaB => P(9)(105),lamdaOut => P(8)(104));
G9105: entity G port map(lamdaA => P(9)(104),lamdaB => P(9)(105),s => s(9)(52),lamdaOut => P(8)(105));
F9106: entity F port map(lamdaA => P(9)(106),lamdaB => P(9)(107),lamdaOut => P(8)(106));
G9107: entity G port map(lamdaA => P(9)(106),lamdaB => P(9)(107),s => s(9)(53),lamdaOut => P(8)(107));
F9108: entity F port map(lamdaA => P(9)(108),lamdaB => P(9)(109),lamdaOut => P(8)(108));
G9109: entity G port map(lamdaA => P(9)(108),lamdaB => P(9)(109),s => s(9)(54),lamdaOut => P(8)(109));
F9110: entity F port map(lamdaA => P(9)(110),lamdaB => P(9)(111),lamdaOut => P(8)(110));
G9111: entity G port map(lamdaA => P(9)(110),lamdaB => P(9)(111),s => s(9)(55),lamdaOut => P(8)(111));
F9112: entity F port map(lamdaA => P(9)(112),lamdaB => P(9)(113),lamdaOut => P(8)(112));
G9113: entity G port map(lamdaA => P(9)(112),lamdaB => P(9)(113),s => s(9)(56),lamdaOut => P(8)(113));
F9114: entity F port map(lamdaA => P(9)(114),lamdaB => P(9)(115),lamdaOut => P(8)(114));
G9115: entity G port map(lamdaA => P(9)(114),lamdaB => P(9)(115),s => s(9)(57),lamdaOut => P(8)(115));
F9116: entity F port map(lamdaA => P(9)(116),lamdaB => P(9)(117),lamdaOut => P(8)(116));
G9117: entity G port map(lamdaA => P(9)(116),lamdaB => P(9)(117),s => s(9)(58),lamdaOut => P(8)(117));
F9118: entity F port map(lamdaA => P(9)(118),lamdaB => P(9)(119),lamdaOut => P(8)(118));
G9119: entity G port map(lamdaA => P(9)(118),lamdaB => P(9)(119),s => s(9)(59),lamdaOut => P(8)(119));
F9120: entity F port map(lamdaA => P(9)(120),lamdaB => P(9)(121),lamdaOut => P(8)(120));
G9121: entity G port map(lamdaA => P(9)(120),lamdaB => P(9)(121),s => s(9)(60),lamdaOut => P(8)(121));
F9122: entity F port map(lamdaA => P(9)(122),lamdaB => P(9)(123),lamdaOut => P(8)(122));
G9123: entity G port map(lamdaA => P(9)(122),lamdaB => P(9)(123),s => s(9)(61),lamdaOut => P(8)(123));
F9124: entity F port map(lamdaA => P(9)(124),lamdaB => P(9)(125),lamdaOut => P(8)(124));
G9125: entity G port map(lamdaA => P(9)(124),lamdaB => P(9)(125),s => s(9)(62),lamdaOut => P(8)(125));
F9126: entity F port map(lamdaA => P(9)(126),lamdaB => P(9)(127),lamdaOut => P(8)(126));
G9127: entity G port map(lamdaA => P(9)(126),lamdaB => P(9)(127),s => s(9)(63),lamdaOut => P(8)(127));
F9128: entity F port map(lamdaA => P(9)(128),lamdaB => P(9)(129),lamdaOut => P(8)(128));
G9129: entity G port map(lamdaA => P(9)(128),lamdaB => P(9)(129),s => s(9)(64),lamdaOut => P(8)(129));
F9130: entity F port map(lamdaA => P(9)(130),lamdaB => P(9)(131),lamdaOut => P(8)(130));
G9131: entity G port map(lamdaA => P(9)(130),lamdaB => P(9)(131),s => s(9)(65),lamdaOut => P(8)(131));
F9132: entity F port map(lamdaA => P(9)(132),lamdaB => P(9)(133),lamdaOut => P(8)(132));
G9133: entity G port map(lamdaA => P(9)(132),lamdaB => P(9)(133),s => s(9)(66),lamdaOut => P(8)(133));
F9134: entity F port map(lamdaA => P(9)(134),lamdaB => P(9)(135),lamdaOut => P(8)(134));
G9135: entity G port map(lamdaA => P(9)(134),lamdaB => P(9)(135),s => s(9)(67),lamdaOut => P(8)(135));
F9136: entity F port map(lamdaA => P(9)(136),lamdaB => P(9)(137),lamdaOut => P(8)(136));
G9137: entity G port map(lamdaA => P(9)(136),lamdaB => P(9)(137),s => s(9)(68),lamdaOut => P(8)(137));
F9138: entity F port map(lamdaA => P(9)(138),lamdaB => P(9)(139),lamdaOut => P(8)(138));
G9139: entity G port map(lamdaA => P(9)(138),lamdaB => P(9)(139),s => s(9)(69),lamdaOut => P(8)(139));
F9140: entity F port map(lamdaA => P(9)(140),lamdaB => P(9)(141),lamdaOut => P(8)(140));
G9141: entity G port map(lamdaA => P(9)(140),lamdaB => P(9)(141),s => s(9)(70),lamdaOut => P(8)(141));
F9142: entity F port map(lamdaA => P(9)(142),lamdaB => P(9)(143),lamdaOut => P(8)(142));
G9143: entity G port map(lamdaA => P(9)(142),lamdaB => P(9)(143),s => s(9)(71),lamdaOut => P(8)(143));
F9144: entity F port map(lamdaA => P(9)(144),lamdaB => P(9)(145),lamdaOut => P(8)(144));
G9145: entity G port map(lamdaA => P(9)(144),lamdaB => P(9)(145),s => s(9)(72),lamdaOut => P(8)(145));
F9146: entity F port map(lamdaA => P(9)(146),lamdaB => P(9)(147),lamdaOut => P(8)(146));
G9147: entity G port map(lamdaA => P(9)(146),lamdaB => P(9)(147),s => s(9)(73),lamdaOut => P(8)(147));
F9148: entity F port map(lamdaA => P(9)(148),lamdaB => P(9)(149),lamdaOut => P(8)(148));
G9149: entity G port map(lamdaA => P(9)(148),lamdaB => P(9)(149),s => s(9)(74),lamdaOut => P(8)(149));
F9150: entity F port map(lamdaA => P(9)(150),lamdaB => P(9)(151),lamdaOut => P(8)(150));
G9151: entity G port map(lamdaA => P(9)(150),lamdaB => P(9)(151),s => s(9)(75),lamdaOut => P(8)(151));
F9152: entity F port map(lamdaA => P(9)(152),lamdaB => P(9)(153),lamdaOut => P(8)(152));
G9153: entity G port map(lamdaA => P(9)(152),lamdaB => P(9)(153),s => s(9)(76),lamdaOut => P(8)(153));
F9154: entity F port map(lamdaA => P(9)(154),lamdaB => P(9)(155),lamdaOut => P(8)(154));
G9155: entity G port map(lamdaA => P(9)(154),lamdaB => P(9)(155),s => s(9)(77),lamdaOut => P(8)(155));
F9156: entity F port map(lamdaA => P(9)(156),lamdaB => P(9)(157),lamdaOut => P(8)(156));
G9157: entity G port map(lamdaA => P(9)(156),lamdaB => P(9)(157),s => s(9)(78),lamdaOut => P(8)(157));
F9158: entity F port map(lamdaA => P(9)(158),lamdaB => P(9)(159),lamdaOut => P(8)(158));
G9159: entity G port map(lamdaA => P(9)(158),lamdaB => P(9)(159),s => s(9)(79),lamdaOut => P(8)(159));
F9160: entity F port map(lamdaA => P(9)(160),lamdaB => P(9)(161),lamdaOut => P(8)(160));
G9161: entity G port map(lamdaA => P(9)(160),lamdaB => P(9)(161),s => s(9)(80),lamdaOut => P(8)(161));
F9162: entity F port map(lamdaA => P(9)(162),lamdaB => P(9)(163),lamdaOut => P(8)(162));
G9163: entity G port map(lamdaA => P(9)(162),lamdaB => P(9)(163),s => s(9)(81),lamdaOut => P(8)(163));
F9164: entity F port map(lamdaA => P(9)(164),lamdaB => P(9)(165),lamdaOut => P(8)(164));
G9165: entity G port map(lamdaA => P(9)(164),lamdaB => P(9)(165),s => s(9)(82),lamdaOut => P(8)(165));
F9166: entity F port map(lamdaA => P(9)(166),lamdaB => P(9)(167),lamdaOut => P(8)(166));
G9167: entity G port map(lamdaA => P(9)(166),lamdaB => P(9)(167),s => s(9)(83),lamdaOut => P(8)(167));
F9168: entity F port map(lamdaA => P(9)(168),lamdaB => P(9)(169),lamdaOut => P(8)(168));
G9169: entity G port map(lamdaA => P(9)(168),lamdaB => P(9)(169),s => s(9)(84),lamdaOut => P(8)(169));
F9170: entity F port map(lamdaA => P(9)(170),lamdaB => P(9)(171),lamdaOut => P(8)(170));
G9171: entity G port map(lamdaA => P(9)(170),lamdaB => P(9)(171),s => s(9)(85),lamdaOut => P(8)(171));
F9172: entity F port map(lamdaA => P(9)(172),lamdaB => P(9)(173),lamdaOut => P(8)(172));
G9173: entity G port map(lamdaA => P(9)(172),lamdaB => P(9)(173),s => s(9)(86),lamdaOut => P(8)(173));
F9174: entity F port map(lamdaA => P(9)(174),lamdaB => P(9)(175),lamdaOut => P(8)(174));
G9175: entity G port map(lamdaA => P(9)(174),lamdaB => P(9)(175),s => s(9)(87),lamdaOut => P(8)(175));
F9176: entity F port map(lamdaA => P(9)(176),lamdaB => P(9)(177),lamdaOut => P(8)(176));
G9177: entity G port map(lamdaA => P(9)(176),lamdaB => P(9)(177),s => s(9)(88),lamdaOut => P(8)(177));
F9178: entity F port map(lamdaA => P(9)(178),lamdaB => P(9)(179),lamdaOut => P(8)(178));
G9179: entity G port map(lamdaA => P(9)(178),lamdaB => P(9)(179),s => s(9)(89),lamdaOut => P(8)(179));
F9180: entity F port map(lamdaA => P(9)(180),lamdaB => P(9)(181),lamdaOut => P(8)(180));
G9181: entity G port map(lamdaA => P(9)(180),lamdaB => P(9)(181),s => s(9)(90),lamdaOut => P(8)(181));
F9182: entity F port map(lamdaA => P(9)(182),lamdaB => P(9)(183),lamdaOut => P(8)(182));
G9183: entity G port map(lamdaA => P(9)(182),lamdaB => P(9)(183),s => s(9)(91),lamdaOut => P(8)(183));
F9184: entity F port map(lamdaA => P(9)(184),lamdaB => P(9)(185),lamdaOut => P(8)(184));
G9185: entity G port map(lamdaA => P(9)(184),lamdaB => P(9)(185),s => s(9)(92),lamdaOut => P(8)(185));
F9186: entity F port map(lamdaA => P(9)(186),lamdaB => P(9)(187),lamdaOut => P(8)(186));
G9187: entity G port map(lamdaA => P(9)(186),lamdaB => P(9)(187),s => s(9)(93),lamdaOut => P(8)(187));
F9188: entity F port map(lamdaA => P(9)(188),lamdaB => P(9)(189),lamdaOut => P(8)(188));
G9189: entity G port map(lamdaA => P(9)(188),lamdaB => P(9)(189),s => s(9)(94),lamdaOut => P(8)(189));
F9190: entity F port map(lamdaA => P(9)(190),lamdaB => P(9)(191),lamdaOut => P(8)(190));
G9191: entity G port map(lamdaA => P(9)(190),lamdaB => P(9)(191),s => s(9)(95),lamdaOut => P(8)(191));
F9192: entity F port map(lamdaA => P(9)(192),lamdaB => P(9)(193),lamdaOut => P(8)(192));
G9193: entity G port map(lamdaA => P(9)(192),lamdaB => P(9)(193),s => s(9)(96),lamdaOut => P(8)(193));
F9194: entity F port map(lamdaA => P(9)(194),lamdaB => P(9)(195),lamdaOut => P(8)(194));
G9195: entity G port map(lamdaA => P(9)(194),lamdaB => P(9)(195),s => s(9)(97),lamdaOut => P(8)(195));
F9196: entity F port map(lamdaA => P(9)(196),lamdaB => P(9)(197),lamdaOut => P(8)(196));
G9197: entity G port map(lamdaA => P(9)(196),lamdaB => P(9)(197),s => s(9)(98),lamdaOut => P(8)(197));
F9198: entity F port map(lamdaA => P(9)(198),lamdaB => P(9)(199),lamdaOut => P(8)(198));
G9199: entity G port map(lamdaA => P(9)(198),lamdaB => P(9)(199),s => s(9)(99),lamdaOut => P(8)(199));
F9200: entity F port map(lamdaA => P(9)(200),lamdaB => P(9)(201),lamdaOut => P(8)(200));
G9201: entity G port map(lamdaA => P(9)(200),lamdaB => P(9)(201),s => s(9)(100),lamdaOut => P(8)(201));
F9202: entity F port map(lamdaA => P(9)(202),lamdaB => P(9)(203),lamdaOut => P(8)(202));
G9203: entity G port map(lamdaA => P(9)(202),lamdaB => P(9)(203),s => s(9)(101),lamdaOut => P(8)(203));
F9204: entity F port map(lamdaA => P(9)(204),lamdaB => P(9)(205),lamdaOut => P(8)(204));
G9205: entity G port map(lamdaA => P(9)(204),lamdaB => P(9)(205),s => s(9)(102),lamdaOut => P(8)(205));
F9206: entity F port map(lamdaA => P(9)(206),lamdaB => P(9)(207),lamdaOut => P(8)(206));
G9207: entity G port map(lamdaA => P(9)(206),lamdaB => P(9)(207),s => s(9)(103),lamdaOut => P(8)(207));
F9208: entity F port map(lamdaA => P(9)(208),lamdaB => P(9)(209),lamdaOut => P(8)(208));
G9209: entity G port map(lamdaA => P(9)(208),lamdaB => P(9)(209),s => s(9)(104),lamdaOut => P(8)(209));
F9210: entity F port map(lamdaA => P(9)(210),lamdaB => P(9)(211),lamdaOut => P(8)(210));
G9211: entity G port map(lamdaA => P(9)(210),lamdaB => P(9)(211),s => s(9)(105),lamdaOut => P(8)(211));
F9212: entity F port map(lamdaA => P(9)(212),lamdaB => P(9)(213),lamdaOut => P(8)(212));
G9213: entity G port map(lamdaA => P(9)(212),lamdaB => P(9)(213),s => s(9)(106),lamdaOut => P(8)(213));
F9214: entity F port map(lamdaA => P(9)(214),lamdaB => P(9)(215),lamdaOut => P(8)(214));
G9215: entity G port map(lamdaA => P(9)(214),lamdaB => P(9)(215),s => s(9)(107),lamdaOut => P(8)(215));
F9216: entity F port map(lamdaA => P(9)(216),lamdaB => P(9)(217),lamdaOut => P(8)(216));
G9217: entity G port map(lamdaA => P(9)(216),lamdaB => P(9)(217),s => s(9)(108),lamdaOut => P(8)(217));
F9218: entity F port map(lamdaA => P(9)(218),lamdaB => P(9)(219),lamdaOut => P(8)(218));
G9219: entity G port map(lamdaA => P(9)(218),lamdaB => P(9)(219),s => s(9)(109),lamdaOut => P(8)(219));
F9220: entity F port map(lamdaA => P(9)(220),lamdaB => P(9)(221),lamdaOut => P(8)(220));
G9221: entity G port map(lamdaA => P(9)(220),lamdaB => P(9)(221),s => s(9)(110),lamdaOut => P(8)(221));
F9222: entity F port map(lamdaA => P(9)(222),lamdaB => P(9)(223),lamdaOut => P(8)(222));
G9223: entity G port map(lamdaA => P(9)(222),lamdaB => P(9)(223),s => s(9)(111),lamdaOut => P(8)(223));
F9224: entity F port map(lamdaA => P(9)(224),lamdaB => P(9)(225),lamdaOut => P(8)(224));
G9225: entity G port map(lamdaA => P(9)(224),lamdaB => P(9)(225),s => s(9)(112),lamdaOut => P(8)(225));
F9226: entity F port map(lamdaA => P(9)(226),lamdaB => P(9)(227),lamdaOut => P(8)(226));
G9227: entity G port map(lamdaA => P(9)(226),lamdaB => P(9)(227),s => s(9)(113),lamdaOut => P(8)(227));
F9228: entity F port map(lamdaA => P(9)(228),lamdaB => P(9)(229),lamdaOut => P(8)(228));
G9229: entity G port map(lamdaA => P(9)(228),lamdaB => P(9)(229),s => s(9)(114),lamdaOut => P(8)(229));
F9230: entity F port map(lamdaA => P(9)(230),lamdaB => P(9)(231),lamdaOut => P(8)(230));
G9231: entity G port map(lamdaA => P(9)(230),lamdaB => P(9)(231),s => s(9)(115),lamdaOut => P(8)(231));
F9232: entity F port map(lamdaA => P(9)(232),lamdaB => P(9)(233),lamdaOut => P(8)(232));
G9233: entity G port map(lamdaA => P(9)(232),lamdaB => P(9)(233),s => s(9)(116),lamdaOut => P(8)(233));
F9234: entity F port map(lamdaA => P(9)(234),lamdaB => P(9)(235),lamdaOut => P(8)(234));
G9235: entity G port map(lamdaA => P(9)(234),lamdaB => P(9)(235),s => s(9)(117),lamdaOut => P(8)(235));
F9236: entity F port map(lamdaA => P(9)(236),lamdaB => P(9)(237),lamdaOut => P(8)(236));
G9237: entity G port map(lamdaA => P(9)(236),lamdaB => P(9)(237),s => s(9)(118),lamdaOut => P(8)(237));
F9238: entity F port map(lamdaA => P(9)(238),lamdaB => P(9)(239),lamdaOut => P(8)(238));
G9239: entity G port map(lamdaA => P(9)(238),lamdaB => P(9)(239),s => s(9)(119),lamdaOut => P(8)(239));
F9240: entity F port map(lamdaA => P(9)(240),lamdaB => P(9)(241),lamdaOut => P(8)(240));
G9241: entity G port map(lamdaA => P(9)(240),lamdaB => P(9)(241),s => s(9)(120),lamdaOut => P(8)(241));
F9242: entity F port map(lamdaA => P(9)(242),lamdaB => P(9)(243),lamdaOut => P(8)(242));
G9243: entity G port map(lamdaA => P(9)(242),lamdaB => P(9)(243),s => s(9)(121),lamdaOut => P(8)(243));
F9244: entity F port map(lamdaA => P(9)(244),lamdaB => P(9)(245),lamdaOut => P(8)(244));
G9245: entity G port map(lamdaA => P(9)(244),lamdaB => P(9)(245),s => s(9)(122),lamdaOut => P(8)(245));
F9246: entity F port map(lamdaA => P(9)(246),lamdaB => P(9)(247),lamdaOut => P(8)(246));
G9247: entity G port map(lamdaA => P(9)(246),lamdaB => P(9)(247),s => s(9)(123),lamdaOut => P(8)(247));
F9248: entity F port map(lamdaA => P(9)(248),lamdaB => P(9)(249),lamdaOut => P(8)(248));
G9249: entity G port map(lamdaA => P(9)(248),lamdaB => P(9)(249),s => s(9)(124),lamdaOut => P(8)(249));
F9250: entity F port map(lamdaA => P(9)(250),lamdaB => P(9)(251),lamdaOut => P(8)(250));
G9251: entity G port map(lamdaA => P(9)(250),lamdaB => P(9)(251),s => s(9)(125),lamdaOut => P(8)(251));
F9252: entity F port map(lamdaA => P(9)(252),lamdaB => P(9)(253),lamdaOut => P(8)(252));
G9253: entity G port map(lamdaA => P(9)(252),lamdaB => P(9)(253),s => s(9)(126),lamdaOut => P(8)(253));
F9254: entity F port map(lamdaA => P(9)(254),lamdaB => P(9)(255),lamdaOut => P(8)(254));
G9255: entity G port map(lamdaA => P(9)(254),lamdaB => P(9)(255),s => s(9)(127),lamdaOut => P(8)(255));
F9256: entity F port map(lamdaA => P(9)(256),lamdaB => P(9)(257),lamdaOut => P(8)(256));
G9257: entity G port map(lamdaA => P(9)(256),lamdaB => P(9)(257),s => s(9)(128),lamdaOut => P(8)(257));
F9258: entity F port map(lamdaA => P(9)(258),lamdaB => P(9)(259),lamdaOut => P(8)(258));
G9259: entity G port map(lamdaA => P(9)(258),lamdaB => P(9)(259),s => s(9)(129),lamdaOut => P(8)(259));
F9260: entity F port map(lamdaA => P(9)(260),lamdaB => P(9)(261),lamdaOut => P(8)(260));
G9261: entity G port map(lamdaA => P(9)(260),lamdaB => P(9)(261),s => s(9)(130),lamdaOut => P(8)(261));
F9262: entity F port map(lamdaA => P(9)(262),lamdaB => P(9)(263),lamdaOut => P(8)(262));
G9263: entity G port map(lamdaA => P(9)(262),lamdaB => P(9)(263),s => s(9)(131),lamdaOut => P(8)(263));
F9264: entity F port map(lamdaA => P(9)(264),lamdaB => P(9)(265),lamdaOut => P(8)(264));
G9265: entity G port map(lamdaA => P(9)(264),lamdaB => P(9)(265),s => s(9)(132),lamdaOut => P(8)(265));
F9266: entity F port map(lamdaA => P(9)(266),lamdaB => P(9)(267),lamdaOut => P(8)(266));
G9267: entity G port map(lamdaA => P(9)(266),lamdaB => P(9)(267),s => s(9)(133),lamdaOut => P(8)(267));
F9268: entity F port map(lamdaA => P(9)(268),lamdaB => P(9)(269),lamdaOut => P(8)(268));
G9269: entity G port map(lamdaA => P(9)(268),lamdaB => P(9)(269),s => s(9)(134),lamdaOut => P(8)(269));
F9270: entity F port map(lamdaA => P(9)(270),lamdaB => P(9)(271),lamdaOut => P(8)(270));
G9271: entity G port map(lamdaA => P(9)(270),lamdaB => P(9)(271),s => s(9)(135),lamdaOut => P(8)(271));
F9272: entity F port map(lamdaA => P(9)(272),lamdaB => P(9)(273),lamdaOut => P(8)(272));
G9273: entity G port map(lamdaA => P(9)(272),lamdaB => P(9)(273),s => s(9)(136),lamdaOut => P(8)(273));
F9274: entity F port map(lamdaA => P(9)(274),lamdaB => P(9)(275),lamdaOut => P(8)(274));
G9275: entity G port map(lamdaA => P(9)(274),lamdaB => P(9)(275),s => s(9)(137),lamdaOut => P(8)(275));
F9276: entity F port map(lamdaA => P(9)(276),lamdaB => P(9)(277),lamdaOut => P(8)(276));
G9277: entity G port map(lamdaA => P(9)(276),lamdaB => P(9)(277),s => s(9)(138),lamdaOut => P(8)(277));
F9278: entity F port map(lamdaA => P(9)(278),lamdaB => P(9)(279),lamdaOut => P(8)(278));
G9279: entity G port map(lamdaA => P(9)(278),lamdaB => P(9)(279),s => s(9)(139),lamdaOut => P(8)(279));
F9280: entity F port map(lamdaA => P(9)(280),lamdaB => P(9)(281),lamdaOut => P(8)(280));
G9281: entity G port map(lamdaA => P(9)(280),lamdaB => P(9)(281),s => s(9)(140),lamdaOut => P(8)(281));
F9282: entity F port map(lamdaA => P(9)(282),lamdaB => P(9)(283),lamdaOut => P(8)(282));
G9283: entity G port map(lamdaA => P(9)(282),lamdaB => P(9)(283),s => s(9)(141),lamdaOut => P(8)(283));
F9284: entity F port map(lamdaA => P(9)(284),lamdaB => P(9)(285),lamdaOut => P(8)(284));
G9285: entity G port map(lamdaA => P(9)(284),lamdaB => P(9)(285),s => s(9)(142),lamdaOut => P(8)(285));
F9286: entity F port map(lamdaA => P(9)(286),lamdaB => P(9)(287),lamdaOut => P(8)(286));
G9287: entity G port map(lamdaA => P(9)(286),lamdaB => P(9)(287),s => s(9)(143),lamdaOut => P(8)(287));
F9288: entity F port map(lamdaA => P(9)(288),lamdaB => P(9)(289),lamdaOut => P(8)(288));
G9289: entity G port map(lamdaA => P(9)(288),lamdaB => P(9)(289),s => s(9)(144),lamdaOut => P(8)(289));
F9290: entity F port map(lamdaA => P(9)(290),lamdaB => P(9)(291),lamdaOut => P(8)(290));
G9291: entity G port map(lamdaA => P(9)(290),lamdaB => P(9)(291),s => s(9)(145),lamdaOut => P(8)(291));
F9292: entity F port map(lamdaA => P(9)(292),lamdaB => P(9)(293),lamdaOut => P(8)(292));
G9293: entity G port map(lamdaA => P(9)(292),lamdaB => P(9)(293),s => s(9)(146),lamdaOut => P(8)(293));
F9294: entity F port map(lamdaA => P(9)(294),lamdaB => P(9)(295),lamdaOut => P(8)(294));
G9295: entity G port map(lamdaA => P(9)(294),lamdaB => P(9)(295),s => s(9)(147),lamdaOut => P(8)(295));
F9296: entity F port map(lamdaA => P(9)(296),lamdaB => P(9)(297),lamdaOut => P(8)(296));
G9297: entity G port map(lamdaA => P(9)(296),lamdaB => P(9)(297),s => s(9)(148),lamdaOut => P(8)(297));
F9298: entity F port map(lamdaA => P(9)(298),lamdaB => P(9)(299),lamdaOut => P(8)(298));
G9299: entity G port map(lamdaA => P(9)(298),lamdaB => P(9)(299),s => s(9)(149),lamdaOut => P(8)(299));
F9300: entity F port map(lamdaA => P(9)(300),lamdaB => P(9)(301),lamdaOut => P(8)(300));
G9301: entity G port map(lamdaA => P(9)(300),lamdaB => P(9)(301),s => s(9)(150),lamdaOut => P(8)(301));
F9302: entity F port map(lamdaA => P(9)(302),lamdaB => P(9)(303),lamdaOut => P(8)(302));
G9303: entity G port map(lamdaA => P(9)(302),lamdaB => P(9)(303),s => s(9)(151),lamdaOut => P(8)(303));
F9304: entity F port map(lamdaA => P(9)(304),lamdaB => P(9)(305),lamdaOut => P(8)(304));
G9305: entity G port map(lamdaA => P(9)(304),lamdaB => P(9)(305),s => s(9)(152),lamdaOut => P(8)(305));
F9306: entity F port map(lamdaA => P(9)(306),lamdaB => P(9)(307),lamdaOut => P(8)(306));
G9307: entity G port map(lamdaA => P(9)(306),lamdaB => P(9)(307),s => s(9)(153),lamdaOut => P(8)(307));
F9308: entity F port map(lamdaA => P(9)(308),lamdaB => P(9)(309),lamdaOut => P(8)(308));
G9309: entity G port map(lamdaA => P(9)(308),lamdaB => P(9)(309),s => s(9)(154),lamdaOut => P(8)(309));
F9310: entity F port map(lamdaA => P(9)(310),lamdaB => P(9)(311),lamdaOut => P(8)(310));
G9311: entity G port map(lamdaA => P(9)(310),lamdaB => P(9)(311),s => s(9)(155),lamdaOut => P(8)(311));
F9312: entity F port map(lamdaA => P(9)(312),lamdaB => P(9)(313),lamdaOut => P(8)(312));
G9313: entity G port map(lamdaA => P(9)(312),lamdaB => P(9)(313),s => s(9)(156),lamdaOut => P(8)(313));
F9314: entity F port map(lamdaA => P(9)(314),lamdaB => P(9)(315),lamdaOut => P(8)(314));
G9315: entity G port map(lamdaA => P(9)(314),lamdaB => P(9)(315),s => s(9)(157),lamdaOut => P(8)(315));
F9316: entity F port map(lamdaA => P(9)(316),lamdaB => P(9)(317),lamdaOut => P(8)(316));
G9317: entity G port map(lamdaA => P(9)(316),lamdaB => P(9)(317),s => s(9)(158),lamdaOut => P(8)(317));
F9318: entity F port map(lamdaA => P(9)(318),lamdaB => P(9)(319),lamdaOut => P(8)(318));
G9319: entity G port map(lamdaA => P(9)(318),lamdaB => P(9)(319),s => s(9)(159),lamdaOut => P(8)(319));
F9320: entity F port map(lamdaA => P(9)(320),lamdaB => P(9)(321),lamdaOut => P(8)(320));
G9321: entity G port map(lamdaA => P(9)(320),lamdaB => P(9)(321),s => s(9)(160),lamdaOut => P(8)(321));
F9322: entity F port map(lamdaA => P(9)(322),lamdaB => P(9)(323),lamdaOut => P(8)(322));
G9323: entity G port map(lamdaA => P(9)(322),lamdaB => P(9)(323),s => s(9)(161),lamdaOut => P(8)(323));
F9324: entity F port map(lamdaA => P(9)(324),lamdaB => P(9)(325),lamdaOut => P(8)(324));
G9325: entity G port map(lamdaA => P(9)(324),lamdaB => P(9)(325),s => s(9)(162),lamdaOut => P(8)(325));
F9326: entity F port map(lamdaA => P(9)(326),lamdaB => P(9)(327),lamdaOut => P(8)(326));
G9327: entity G port map(lamdaA => P(9)(326),lamdaB => P(9)(327),s => s(9)(163),lamdaOut => P(8)(327));
F9328: entity F port map(lamdaA => P(9)(328),lamdaB => P(9)(329),lamdaOut => P(8)(328));
G9329: entity G port map(lamdaA => P(9)(328),lamdaB => P(9)(329),s => s(9)(164),lamdaOut => P(8)(329));
F9330: entity F port map(lamdaA => P(9)(330),lamdaB => P(9)(331),lamdaOut => P(8)(330));
G9331: entity G port map(lamdaA => P(9)(330),lamdaB => P(9)(331),s => s(9)(165),lamdaOut => P(8)(331));
F9332: entity F port map(lamdaA => P(9)(332),lamdaB => P(9)(333),lamdaOut => P(8)(332));
G9333: entity G port map(lamdaA => P(9)(332),lamdaB => P(9)(333),s => s(9)(166),lamdaOut => P(8)(333));
F9334: entity F port map(lamdaA => P(9)(334),lamdaB => P(9)(335),lamdaOut => P(8)(334));
G9335: entity G port map(lamdaA => P(9)(334),lamdaB => P(9)(335),s => s(9)(167),lamdaOut => P(8)(335));
F9336: entity F port map(lamdaA => P(9)(336),lamdaB => P(9)(337),lamdaOut => P(8)(336));
G9337: entity G port map(lamdaA => P(9)(336),lamdaB => P(9)(337),s => s(9)(168),lamdaOut => P(8)(337));
F9338: entity F port map(lamdaA => P(9)(338),lamdaB => P(9)(339),lamdaOut => P(8)(338));
G9339: entity G port map(lamdaA => P(9)(338),lamdaB => P(9)(339),s => s(9)(169),lamdaOut => P(8)(339));
F9340: entity F port map(lamdaA => P(9)(340),lamdaB => P(9)(341),lamdaOut => P(8)(340));
G9341: entity G port map(lamdaA => P(9)(340),lamdaB => P(9)(341),s => s(9)(170),lamdaOut => P(8)(341));
F9342: entity F port map(lamdaA => P(9)(342),lamdaB => P(9)(343),lamdaOut => P(8)(342));
G9343: entity G port map(lamdaA => P(9)(342),lamdaB => P(9)(343),s => s(9)(171),lamdaOut => P(8)(343));
F9344: entity F port map(lamdaA => P(9)(344),lamdaB => P(9)(345),lamdaOut => P(8)(344));
G9345: entity G port map(lamdaA => P(9)(344),lamdaB => P(9)(345),s => s(9)(172),lamdaOut => P(8)(345));
F9346: entity F port map(lamdaA => P(9)(346),lamdaB => P(9)(347),lamdaOut => P(8)(346));
G9347: entity G port map(lamdaA => P(9)(346),lamdaB => P(9)(347),s => s(9)(173),lamdaOut => P(8)(347));
F9348: entity F port map(lamdaA => P(9)(348),lamdaB => P(9)(349),lamdaOut => P(8)(348));
G9349: entity G port map(lamdaA => P(9)(348),lamdaB => P(9)(349),s => s(9)(174),lamdaOut => P(8)(349));
F9350: entity F port map(lamdaA => P(9)(350),lamdaB => P(9)(351),lamdaOut => P(8)(350));
G9351: entity G port map(lamdaA => P(9)(350),lamdaB => P(9)(351),s => s(9)(175),lamdaOut => P(8)(351));
F9352: entity F port map(lamdaA => P(9)(352),lamdaB => P(9)(353),lamdaOut => P(8)(352));
G9353: entity G port map(lamdaA => P(9)(352),lamdaB => P(9)(353),s => s(9)(176),lamdaOut => P(8)(353));
F9354: entity F port map(lamdaA => P(9)(354),lamdaB => P(9)(355),lamdaOut => P(8)(354));
G9355: entity G port map(lamdaA => P(9)(354),lamdaB => P(9)(355),s => s(9)(177),lamdaOut => P(8)(355));
F9356: entity F port map(lamdaA => P(9)(356),lamdaB => P(9)(357),lamdaOut => P(8)(356));
G9357: entity G port map(lamdaA => P(9)(356),lamdaB => P(9)(357),s => s(9)(178),lamdaOut => P(8)(357));
F9358: entity F port map(lamdaA => P(9)(358),lamdaB => P(9)(359),lamdaOut => P(8)(358));
G9359: entity G port map(lamdaA => P(9)(358),lamdaB => P(9)(359),s => s(9)(179),lamdaOut => P(8)(359));
F9360: entity F port map(lamdaA => P(9)(360),lamdaB => P(9)(361),lamdaOut => P(8)(360));
G9361: entity G port map(lamdaA => P(9)(360),lamdaB => P(9)(361),s => s(9)(180),lamdaOut => P(8)(361));
F9362: entity F port map(lamdaA => P(9)(362),lamdaB => P(9)(363),lamdaOut => P(8)(362));
G9363: entity G port map(lamdaA => P(9)(362),lamdaB => P(9)(363),s => s(9)(181),lamdaOut => P(8)(363));
F9364: entity F port map(lamdaA => P(9)(364),lamdaB => P(9)(365),lamdaOut => P(8)(364));
G9365: entity G port map(lamdaA => P(9)(364),lamdaB => P(9)(365),s => s(9)(182),lamdaOut => P(8)(365));
F9366: entity F port map(lamdaA => P(9)(366),lamdaB => P(9)(367),lamdaOut => P(8)(366));
G9367: entity G port map(lamdaA => P(9)(366),lamdaB => P(9)(367),s => s(9)(183),lamdaOut => P(8)(367));
F9368: entity F port map(lamdaA => P(9)(368),lamdaB => P(9)(369),lamdaOut => P(8)(368));
G9369: entity G port map(lamdaA => P(9)(368),lamdaB => P(9)(369),s => s(9)(184),lamdaOut => P(8)(369));
F9370: entity F port map(lamdaA => P(9)(370),lamdaB => P(9)(371),lamdaOut => P(8)(370));
G9371: entity G port map(lamdaA => P(9)(370),lamdaB => P(9)(371),s => s(9)(185),lamdaOut => P(8)(371));
F9372: entity F port map(lamdaA => P(9)(372),lamdaB => P(9)(373),lamdaOut => P(8)(372));
G9373: entity G port map(lamdaA => P(9)(372),lamdaB => P(9)(373),s => s(9)(186),lamdaOut => P(8)(373));
F9374: entity F port map(lamdaA => P(9)(374),lamdaB => P(9)(375),lamdaOut => P(8)(374));
G9375: entity G port map(lamdaA => P(9)(374),lamdaB => P(9)(375),s => s(9)(187),lamdaOut => P(8)(375));
F9376: entity F port map(lamdaA => P(9)(376),lamdaB => P(9)(377),lamdaOut => P(8)(376));
G9377: entity G port map(lamdaA => P(9)(376),lamdaB => P(9)(377),s => s(9)(188),lamdaOut => P(8)(377));
F9378: entity F port map(lamdaA => P(9)(378),lamdaB => P(9)(379),lamdaOut => P(8)(378));
G9379: entity G port map(lamdaA => P(9)(378),lamdaB => P(9)(379),s => s(9)(189),lamdaOut => P(8)(379));
F9380: entity F port map(lamdaA => P(9)(380),lamdaB => P(9)(381),lamdaOut => P(8)(380));
G9381: entity G port map(lamdaA => P(9)(380),lamdaB => P(9)(381),s => s(9)(190),lamdaOut => P(8)(381));
F9382: entity F port map(lamdaA => P(9)(382),lamdaB => P(9)(383),lamdaOut => P(8)(382));
G9383: entity G port map(lamdaA => P(9)(382),lamdaB => P(9)(383),s => s(9)(191),lamdaOut => P(8)(383));
F9384: entity F port map(lamdaA => P(9)(384),lamdaB => P(9)(385),lamdaOut => P(8)(384));
G9385: entity G port map(lamdaA => P(9)(384),lamdaB => P(9)(385),s => s(9)(192),lamdaOut => P(8)(385));
F9386: entity F port map(lamdaA => P(9)(386),lamdaB => P(9)(387),lamdaOut => P(8)(386));
G9387: entity G port map(lamdaA => P(9)(386),lamdaB => P(9)(387),s => s(9)(193),lamdaOut => P(8)(387));
F9388: entity F port map(lamdaA => P(9)(388),lamdaB => P(9)(389),lamdaOut => P(8)(388));
G9389: entity G port map(lamdaA => P(9)(388),lamdaB => P(9)(389),s => s(9)(194),lamdaOut => P(8)(389));
F9390: entity F port map(lamdaA => P(9)(390),lamdaB => P(9)(391),lamdaOut => P(8)(390));
G9391: entity G port map(lamdaA => P(9)(390),lamdaB => P(9)(391),s => s(9)(195),lamdaOut => P(8)(391));
F9392: entity F port map(lamdaA => P(9)(392),lamdaB => P(9)(393),lamdaOut => P(8)(392));
G9393: entity G port map(lamdaA => P(9)(392),lamdaB => P(9)(393),s => s(9)(196),lamdaOut => P(8)(393));
F9394: entity F port map(lamdaA => P(9)(394),lamdaB => P(9)(395),lamdaOut => P(8)(394));
G9395: entity G port map(lamdaA => P(9)(394),lamdaB => P(9)(395),s => s(9)(197),lamdaOut => P(8)(395));
F9396: entity F port map(lamdaA => P(9)(396),lamdaB => P(9)(397),lamdaOut => P(8)(396));
G9397: entity G port map(lamdaA => P(9)(396),lamdaB => P(9)(397),s => s(9)(198),lamdaOut => P(8)(397));
F9398: entity F port map(lamdaA => P(9)(398),lamdaB => P(9)(399),lamdaOut => P(8)(398));
G9399: entity G port map(lamdaA => P(9)(398),lamdaB => P(9)(399),s => s(9)(199),lamdaOut => P(8)(399));
F9400: entity F port map(lamdaA => P(9)(400),lamdaB => P(9)(401),lamdaOut => P(8)(400));
G9401: entity G port map(lamdaA => P(9)(400),lamdaB => P(9)(401),s => s(9)(200),lamdaOut => P(8)(401));
F9402: entity F port map(lamdaA => P(9)(402),lamdaB => P(9)(403),lamdaOut => P(8)(402));
G9403: entity G port map(lamdaA => P(9)(402),lamdaB => P(9)(403),s => s(9)(201),lamdaOut => P(8)(403));
F9404: entity F port map(lamdaA => P(9)(404),lamdaB => P(9)(405),lamdaOut => P(8)(404));
G9405: entity G port map(lamdaA => P(9)(404),lamdaB => P(9)(405),s => s(9)(202),lamdaOut => P(8)(405));
F9406: entity F port map(lamdaA => P(9)(406),lamdaB => P(9)(407),lamdaOut => P(8)(406));
G9407: entity G port map(lamdaA => P(9)(406),lamdaB => P(9)(407),s => s(9)(203),lamdaOut => P(8)(407));
F9408: entity F port map(lamdaA => P(9)(408),lamdaB => P(9)(409),lamdaOut => P(8)(408));
G9409: entity G port map(lamdaA => P(9)(408),lamdaB => P(9)(409),s => s(9)(204),lamdaOut => P(8)(409));
F9410: entity F port map(lamdaA => P(9)(410),lamdaB => P(9)(411),lamdaOut => P(8)(410));
G9411: entity G port map(lamdaA => P(9)(410),lamdaB => P(9)(411),s => s(9)(205),lamdaOut => P(8)(411));
F9412: entity F port map(lamdaA => P(9)(412),lamdaB => P(9)(413),lamdaOut => P(8)(412));
G9413: entity G port map(lamdaA => P(9)(412),lamdaB => P(9)(413),s => s(9)(206),lamdaOut => P(8)(413));
F9414: entity F port map(lamdaA => P(9)(414),lamdaB => P(9)(415),lamdaOut => P(8)(414));
G9415: entity G port map(lamdaA => P(9)(414),lamdaB => P(9)(415),s => s(9)(207),lamdaOut => P(8)(415));
F9416: entity F port map(lamdaA => P(9)(416),lamdaB => P(9)(417),lamdaOut => P(8)(416));
G9417: entity G port map(lamdaA => P(9)(416),lamdaB => P(9)(417),s => s(9)(208),lamdaOut => P(8)(417));
F9418: entity F port map(lamdaA => P(9)(418),lamdaB => P(9)(419),lamdaOut => P(8)(418));
G9419: entity G port map(lamdaA => P(9)(418),lamdaB => P(9)(419),s => s(9)(209),lamdaOut => P(8)(419));
F9420: entity F port map(lamdaA => P(9)(420),lamdaB => P(9)(421),lamdaOut => P(8)(420));
G9421: entity G port map(lamdaA => P(9)(420),lamdaB => P(9)(421),s => s(9)(210),lamdaOut => P(8)(421));
F9422: entity F port map(lamdaA => P(9)(422),lamdaB => P(9)(423),lamdaOut => P(8)(422));
G9423: entity G port map(lamdaA => P(9)(422),lamdaB => P(9)(423),s => s(9)(211),lamdaOut => P(8)(423));
F9424: entity F port map(lamdaA => P(9)(424),lamdaB => P(9)(425),lamdaOut => P(8)(424));
G9425: entity G port map(lamdaA => P(9)(424),lamdaB => P(9)(425),s => s(9)(212),lamdaOut => P(8)(425));
F9426: entity F port map(lamdaA => P(9)(426),lamdaB => P(9)(427),lamdaOut => P(8)(426));
G9427: entity G port map(lamdaA => P(9)(426),lamdaB => P(9)(427),s => s(9)(213),lamdaOut => P(8)(427));
F9428: entity F port map(lamdaA => P(9)(428),lamdaB => P(9)(429),lamdaOut => P(8)(428));
G9429: entity G port map(lamdaA => P(9)(428),lamdaB => P(9)(429),s => s(9)(214),lamdaOut => P(8)(429));
F9430: entity F port map(lamdaA => P(9)(430),lamdaB => P(9)(431),lamdaOut => P(8)(430));
G9431: entity G port map(lamdaA => P(9)(430),lamdaB => P(9)(431),s => s(9)(215),lamdaOut => P(8)(431));
F9432: entity F port map(lamdaA => P(9)(432),lamdaB => P(9)(433),lamdaOut => P(8)(432));
G9433: entity G port map(lamdaA => P(9)(432),lamdaB => P(9)(433),s => s(9)(216),lamdaOut => P(8)(433));
F9434: entity F port map(lamdaA => P(9)(434),lamdaB => P(9)(435),lamdaOut => P(8)(434));
G9435: entity G port map(lamdaA => P(9)(434),lamdaB => P(9)(435),s => s(9)(217),lamdaOut => P(8)(435));
F9436: entity F port map(lamdaA => P(9)(436),lamdaB => P(9)(437),lamdaOut => P(8)(436));
G9437: entity G port map(lamdaA => P(9)(436),lamdaB => P(9)(437),s => s(9)(218),lamdaOut => P(8)(437));
F9438: entity F port map(lamdaA => P(9)(438),lamdaB => P(9)(439),lamdaOut => P(8)(438));
G9439: entity G port map(lamdaA => P(9)(438),lamdaB => P(9)(439),s => s(9)(219),lamdaOut => P(8)(439));
F9440: entity F port map(lamdaA => P(9)(440),lamdaB => P(9)(441),lamdaOut => P(8)(440));
G9441: entity G port map(lamdaA => P(9)(440),lamdaB => P(9)(441),s => s(9)(220),lamdaOut => P(8)(441));
F9442: entity F port map(lamdaA => P(9)(442),lamdaB => P(9)(443),lamdaOut => P(8)(442));
G9443: entity G port map(lamdaA => P(9)(442),lamdaB => P(9)(443),s => s(9)(221),lamdaOut => P(8)(443));
F9444: entity F port map(lamdaA => P(9)(444),lamdaB => P(9)(445),lamdaOut => P(8)(444));
G9445: entity G port map(lamdaA => P(9)(444),lamdaB => P(9)(445),s => s(9)(222),lamdaOut => P(8)(445));
F9446: entity F port map(lamdaA => P(9)(446),lamdaB => P(9)(447),lamdaOut => P(8)(446));
G9447: entity G port map(lamdaA => P(9)(446),lamdaB => P(9)(447),s => s(9)(223),lamdaOut => P(8)(447));
F9448: entity F port map(lamdaA => P(9)(448),lamdaB => P(9)(449),lamdaOut => P(8)(448));
G9449: entity G port map(lamdaA => P(9)(448),lamdaB => P(9)(449),s => s(9)(224),lamdaOut => P(8)(449));
F9450: entity F port map(lamdaA => P(9)(450),lamdaB => P(9)(451),lamdaOut => P(8)(450));
G9451: entity G port map(lamdaA => P(9)(450),lamdaB => P(9)(451),s => s(9)(225),lamdaOut => P(8)(451));
F9452: entity F port map(lamdaA => P(9)(452),lamdaB => P(9)(453),lamdaOut => P(8)(452));
G9453: entity G port map(lamdaA => P(9)(452),lamdaB => P(9)(453),s => s(9)(226),lamdaOut => P(8)(453));
F9454: entity F port map(lamdaA => P(9)(454),lamdaB => P(9)(455),lamdaOut => P(8)(454));
G9455: entity G port map(lamdaA => P(9)(454),lamdaB => P(9)(455),s => s(9)(227),lamdaOut => P(8)(455));
F9456: entity F port map(lamdaA => P(9)(456),lamdaB => P(9)(457),lamdaOut => P(8)(456));
G9457: entity G port map(lamdaA => P(9)(456),lamdaB => P(9)(457),s => s(9)(228),lamdaOut => P(8)(457));
F9458: entity F port map(lamdaA => P(9)(458),lamdaB => P(9)(459),lamdaOut => P(8)(458));
G9459: entity G port map(lamdaA => P(9)(458),lamdaB => P(9)(459),s => s(9)(229),lamdaOut => P(8)(459));
F9460: entity F port map(lamdaA => P(9)(460),lamdaB => P(9)(461),lamdaOut => P(8)(460));
G9461: entity G port map(lamdaA => P(9)(460),lamdaB => P(9)(461),s => s(9)(230),lamdaOut => P(8)(461));
F9462: entity F port map(lamdaA => P(9)(462),lamdaB => P(9)(463),lamdaOut => P(8)(462));
G9463: entity G port map(lamdaA => P(9)(462),lamdaB => P(9)(463),s => s(9)(231),lamdaOut => P(8)(463));
F9464: entity F port map(lamdaA => P(9)(464),lamdaB => P(9)(465),lamdaOut => P(8)(464));
G9465: entity G port map(lamdaA => P(9)(464),lamdaB => P(9)(465),s => s(9)(232),lamdaOut => P(8)(465));
F9466: entity F port map(lamdaA => P(9)(466),lamdaB => P(9)(467),lamdaOut => P(8)(466));
G9467: entity G port map(lamdaA => P(9)(466),lamdaB => P(9)(467),s => s(9)(233),lamdaOut => P(8)(467));
F9468: entity F port map(lamdaA => P(9)(468),lamdaB => P(9)(469),lamdaOut => P(8)(468));
G9469: entity G port map(lamdaA => P(9)(468),lamdaB => P(9)(469),s => s(9)(234),lamdaOut => P(8)(469));
F9470: entity F port map(lamdaA => P(9)(470),lamdaB => P(9)(471),lamdaOut => P(8)(470));
G9471: entity G port map(lamdaA => P(9)(470),lamdaB => P(9)(471),s => s(9)(235),lamdaOut => P(8)(471));
F9472: entity F port map(lamdaA => P(9)(472),lamdaB => P(9)(473),lamdaOut => P(8)(472));
G9473: entity G port map(lamdaA => P(9)(472),lamdaB => P(9)(473),s => s(9)(236),lamdaOut => P(8)(473));
F9474: entity F port map(lamdaA => P(9)(474),lamdaB => P(9)(475),lamdaOut => P(8)(474));
G9475: entity G port map(lamdaA => P(9)(474),lamdaB => P(9)(475),s => s(9)(237),lamdaOut => P(8)(475));
F9476: entity F port map(lamdaA => P(9)(476),lamdaB => P(9)(477),lamdaOut => P(8)(476));
G9477: entity G port map(lamdaA => P(9)(476),lamdaB => P(9)(477),s => s(9)(238),lamdaOut => P(8)(477));
F9478: entity F port map(lamdaA => P(9)(478),lamdaB => P(9)(479),lamdaOut => P(8)(478));
G9479: entity G port map(lamdaA => P(9)(478),lamdaB => P(9)(479),s => s(9)(239),lamdaOut => P(8)(479));
F9480: entity F port map(lamdaA => P(9)(480),lamdaB => P(9)(481),lamdaOut => P(8)(480));
G9481: entity G port map(lamdaA => P(9)(480),lamdaB => P(9)(481),s => s(9)(240),lamdaOut => P(8)(481));
F9482: entity F port map(lamdaA => P(9)(482),lamdaB => P(9)(483),lamdaOut => P(8)(482));
G9483: entity G port map(lamdaA => P(9)(482),lamdaB => P(9)(483),s => s(9)(241),lamdaOut => P(8)(483));
F9484: entity F port map(lamdaA => P(9)(484),lamdaB => P(9)(485),lamdaOut => P(8)(484));
G9485: entity G port map(lamdaA => P(9)(484),lamdaB => P(9)(485),s => s(9)(242),lamdaOut => P(8)(485));
F9486: entity F port map(lamdaA => P(9)(486),lamdaB => P(9)(487),lamdaOut => P(8)(486));
G9487: entity G port map(lamdaA => P(9)(486),lamdaB => P(9)(487),s => s(9)(243),lamdaOut => P(8)(487));
F9488: entity F port map(lamdaA => P(9)(488),lamdaB => P(9)(489),lamdaOut => P(8)(488));
G9489: entity G port map(lamdaA => P(9)(488),lamdaB => P(9)(489),s => s(9)(244),lamdaOut => P(8)(489));
F9490: entity F port map(lamdaA => P(9)(490),lamdaB => P(9)(491),lamdaOut => P(8)(490));
G9491: entity G port map(lamdaA => P(9)(490),lamdaB => P(9)(491),s => s(9)(245),lamdaOut => P(8)(491));
F9492: entity F port map(lamdaA => P(9)(492),lamdaB => P(9)(493),lamdaOut => P(8)(492));
G9493: entity G port map(lamdaA => P(9)(492),lamdaB => P(9)(493),s => s(9)(246),lamdaOut => P(8)(493));
F9494: entity F port map(lamdaA => P(9)(494),lamdaB => P(9)(495),lamdaOut => P(8)(494));
G9495: entity G port map(lamdaA => P(9)(494),lamdaB => P(9)(495),s => s(9)(247),lamdaOut => P(8)(495));
F9496: entity F port map(lamdaA => P(9)(496),lamdaB => P(9)(497),lamdaOut => P(8)(496));
G9497: entity G port map(lamdaA => P(9)(496),lamdaB => P(9)(497),s => s(9)(248),lamdaOut => P(8)(497));
F9498: entity F port map(lamdaA => P(9)(498),lamdaB => P(9)(499),lamdaOut => P(8)(498));
G9499: entity G port map(lamdaA => P(9)(498),lamdaB => P(9)(499),s => s(9)(249),lamdaOut => P(8)(499));
F9500: entity F port map(lamdaA => P(9)(500),lamdaB => P(9)(501),lamdaOut => P(8)(500));
G9501: entity G port map(lamdaA => P(9)(500),lamdaB => P(9)(501),s => s(9)(250),lamdaOut => P(8)(501));
F9502: entity F port map(lamdaA => P(9)(502),lamdaB => P(9)(503),lamdaOut => P(8)(502));
G9503: entity G port map(lamdaA => P(9)(502),lamdaB => P(9)(503),s => s(9)(251),lamdaOut => P(8)(503));
F9504: entity F port map(lamdaA => P(9)(504),lamdaB => P(9)(505),lamdaOut => P(8)(504));
G9505: entity G port map(lamdaA => P(9)(504),lamdaB => P(9)(505),s => s(9)(252),lamdaOut => P(8)(505));
F9506: entity F port map(lamdaA => P(9)(506),lamdaB => P(9)(507),lamdaOut => P(8)(506));
G9507: entity G port map(lamdaA => P(9)(506),lamdaB => P(9)(507),s => s(9)(253),lamdaOut => P(8)(507));
F9508: entity F port map(lamdaA => P(9)(508),lamdaB => P(9)(509),lamdaOut => P(8)(508));
G9509: entity G port map(lamdaA => P(9)(508),lamdaB => P(9)(509),s => s(9)(254),lamdaOut => P(8)(509));
F9510: entity F port map(lamdaA => P(9)(510),lamdaB => P(9)(511),lamdaOut => P(8)(510));
G9511: entity G port map(lamdaA => P(9)(510),lamdaB => P(9)(511),s => s(9)(255),lamdaOut => P(8)(511));
-- STAGE 8
F80: entity F port map(lamdaA => P(8)(0),lamdaB => P(8)(2),lamdaOut => P(7)(0));
F81: entity F port map(lamdaA => P(8)(1),lamdaB => P(8)(3),lamdaOut => P(7)(1));
G82: entity G port map(lamdaA => P(8)(0),lamdaB => P(8)(2),s => s(8)(0),lamdaOut => P(7)(2));
G83: entity G port map(lamdaA => P(8)(1),lamdaB => P(8)(3),s => s(8)(1),lamdaOut => P(7)(3));
F84: entity F port map(lamdaA => P(8)(4),lamdaB => P(8)(6),lamdaOut => P(7)(4));
F85: entity F port map(lamdaA => P(8)(5),lamdaB => P(8)(7),lamdaOut => P(7)(5));
G86: entity G port map(lamdaA => P(8)(4),lamdaB => P(8)(6),s => s(8)(2),lamdaOut => P(7)(6));
G87: entity G port map(lamdaA => P(8)(5),lamdaB => P(8)(7),s => s(8)(3),lamdaOut => P(7)(7));
F88: entity F port map(lamdaA => P(8)(8),lamdaB => P(8)(10),lamdaOut => P(7)(8));
F89: entity F port map(lamdaA => P(8)(9),lamdaB => P(8)(11),lamdaOut => P(7)(9));
G810: entity G port map(lamdaA => P(8)(8),lamdaB => P(8)(10),s => s(8)(4),lamdaOut => P(7)(10));
G811: entity G port map(lamdaA => P(8)(9),lamdaB => P(8)(11),s => s(8)(5),lamdaOut => P(7)(11));
F812: entity F port map(lamdaA => P(8)(12),lamdaB => P(8)(14),lamdaOut => P(7)(12));
F813: entity F port map(lamdaA => P(8)(13),lamdaB => P(8)(15),lamdaOut => P(7)(13));
G814: entity G port map(lamdaA => P(8)(12),lamdaB => P(8)(14),s => s(8)(6),lamdaOut => P(7)(14));
G815: entity G port map(lamdaA => P(8)(13),lamdaB => P(8)(15),s => s(8)(7),lamdaOut => P(7)(15));
F816: entity F port map(lamdaA => P(8)(16),lamdaB => P(8)(18),lamdaOut => P(7)(16));
F817: entity F port map(lamdaA => P(8)(17),lamdaB => P(8)(19),lamdaOut => P(7)(17));
G818: entity G port map(lamdaA => P(8)(16),lamdaB => P(8)(18),s => s(8)(8),lamdaOut => P(7)(18));
G819: entity G port map(lamdaA => P(8)(17),lamdaB => P(8)(19),s => s(8)(9),lamdaOut => P(7)(19));
F820: entity F port map(lamdaA => P(8)(20),lamdaB => P(8)(22),lamdaOut => P(7)(20));
F821: entity F port map(lamdaA => P(8)(21),lamdaB => P(8)(23),lamdaOut => P(7)(21));
G822: entity G port map(lamdaA => P(8)(20),lamdaB => P(8)(22),s => s(8)(10),lamdaOut => P(7)(22));
G823: entity G port map(lamdaA => P(8)(21),lamdaB => P(8)(23),s => s(8)(11),lamdaOut => P(7)(23));
F824: entity F port map(lamdaA => P(8)(24),lamdaB => P(8)(26),lamdaOut => P(7)(24));
F825: entity F port map(lamdaA => P(8)(25),lamdaB => P(8)(27),lamdaOut => P(7)(25));
G826: entity G port map(lamdaA => P(8)(24),lamdaB => P(8)(26),s => s(8)(12),lamdaOut => P(7)(26));
G827: entity G port map(lamdaA => P(8)(25),lamdaB => P(8)(27),s => s(8)(13),lamdaOut => P(7)(27));
F828: entity F port map(lamdaA => P(8)(28),lamdaB => P(8)(30),lamdaOut => P(7)(28));
F829: entity F port map(lamdaA => P(8)(29),lamdaB => P(8)(31),lamdaOut => P(7)(29));
G830: entity G port map(lamdaA => P(8)(28),lamdaB => P(8)(30),s => s(8)(14),lamdaOut => P(7)(30));
G831: entity G port map(lamdaA => P(8)(29),lamdaB => P(8)(31),s => s(8)(15),lamdaOut => P(7)(31));
F832: entity F port map(lamdaA => P(8)(32),lamdaB => P(8)(34),lamdaOut => P(7)(32));
F833: entity F port map(lamdaA => P(8)(33),lamdaB => P(8)(35),lamdaOut => P(7)(33));
G834: entity G port map(lamdaA => P(8)(32),lamdaB => P(8)(34),s => s(8)(16),lamdaOut => P(7)(34));
G835: entity G port map(lamdaA => P(8)(33),lamdaB => P(8)(35),s => s(8)(17),lamdaOut => P(7)(35));
F836: entity F port map(lamdaA => P(8)(36),lamdaB => P(8)(38),lamdaOut => P(7)(36));
F837: entity F port map(lamdaA => P(8)(37),lamdaB => P(8)(39),lamdaOut => P(7)(37));
G838: entity G port map(lamdaA => P(8)(36),lamdaB => P(8)(38),s => s(8)(18),lamdaOut => P(7)(38));
G839: entity G port map(lamdaA => P(8)(37),lamdaB => P(8)(39),s => s(8)(19),lamdaOut => P(7)(39));
F840: entity F port map(lamdaA => P(8)(40),lamdaB => P(8)(42),lamdaOut => P(7)(40));
F841: entity F port map(lamdaA => P(8)(41),lamdaB => P(8)(43),lamdaOut => P(7)(41));
G842: entity G port map(lamdaA => P(8)(40),lamdaB => P(8)(42),s => s(8)(20),lamdaOut => P(7)(42));
G843: entity G port map(lamdaA => P(8)(41),lamdaB => P(8)(43),s => s(8)(21),lamdaOut => P(7)(43));
F844: entity F port map(lamdaA => P(8)(44),lamdaB => P(8)(46),lamdaOut => P(7)(44));
F845: entity F port map(lamdaA => P(8)(45),lamdaB => P(8)(47),lamdaOut => P(7)(45));
G846: entity G port map(lamdaA => P(8)(44),lamdaB => P(8)(46),s => s(8)(22),lamdaOut => P(7)(46));
G847: entity G port map(lamdaA => P(8)(45),lamdaB => P(8)(47),s => s(8)(23),lamdaOut => P(7)(47));
F848: entity F port map(lamdaA => P(8)(48),lamdaB => P(8)(50),lamdaOut => P(7)(48));
F849: entity F port map(lamdaA => P(8)(49),lamdaB => P(8)(51),lamdaOut => P(7)(49));
G850: entity G port map(lamdaA => P(8)(48),lamdaB => P(8)(50),s => s(8)(24),lamdaOut => P(7)(50));
G851: entity G port map(lamdaA => P(8)(49),lamdaB => P(8)(51),s => s(8)(25),lamdaOut => P(7)(51));
F852: entity F port map(lamdaA => P(8)(52),lamdaB => P(8)(54),lamdaOut => P(7)(52));
F853: entity F port map(lamdaA => P(8)(53),lamdaB => P(8)(55),lamdaOut => P(7)(53));
G854: entity G port map(lamdaA => P(8)(52),lamdaB => P(8)(54),s => s(8)(26),lamdaOut => P(7)(54));
G855: entity G port map(lamdaA => P(8)(53),lamdaB => P(8)(55),s => s(8)(27),lamdaOut => P(7)(55));
F856: entity F port map(lamdaA => P(8)(56),lamdaB => P(8)(58),lamdaOut => P(7)(56));
F857: entity F port map(lamdaA => P(8)(57),lamdaB => P(8)(59),lamdaOut => P(7)(57));
G858: entity G port map(lamdaA => P(8)(56),lamdaB => P(8)(58),s => s(8)(28),lamdaOut => P(7)(58));
G859: entity G port map(lamdaA => P(8)(57),lamdaB => P(8)(59),s => s(8)(29),lamdaOut => P(7)(59));
F860: entity F port map(lamdaA => P(8)(60),lamdaB => P(8)(62),lamdaOut => P(7)(60));
F861: entity F port map(lamdaA => P(8)(61),lamdaB => P(8)(63),lamdaOut => P(7)(61));
G862: entity G port map(lamdaA => P(8)(60),lamdaB => P(8)(62),s => s(8)(30),lamdaOut => P(7)(62));
G863: entity G port map(lamdaA => P(8)(61),lamdaB => P(8)(63),s => s(8)(31),lamdaOut => P(7)(63));
F864: entity F port map(lamdaA => P(8)(64),lamdaB => P(8)(66),lamdaOut => P(7)(64));
F865: entity F port map(lamdaA => P(8)(65),lamdaB => P(8)(67),lamdaOut => P(7)(65));
G866: entity G port map(lamdaA => P(8)(64),lamdaB => P(8)(66),s => s(8)(32),lamdaOut => P(7)(66));
G867: entity G port map(lamdaA => P(8)(65),lamdaB => P(8)(67),s => s(8)(33),lamdaOut => P(7)(67));
F868: entity F port map(lamdaA => P(8)(68),lamdaB => P(8)(70),lamdaOut => P(7)(68));
F869: entity F port map(lamdaA => P(8)(69),lamdaB => P(8)(71),lamdaOut => P(7)(69));
G870: entity G port map(lamdaA => P(8)(68),lamdaB => P(8)(70),s => s(8)(34),lamdaOut => P(7)(70));
G871: entity G port map(lamdaA => P(8)(69),lamdaB => P(8)(71),s => s(8)(35),lamdaOut => P(7)(71));
F872: entity F port map(lamdaA => P(8)(72),lamdaB => P(8)(74),lamdaOut => P(7)(72));
F873: entity F port map(lamdaA => P(8)(73),lamdaB => P(8)(75),lamdaOut => P(7)(73));
G874: entity G port map(lamdaA => P(8)(72),lamdaB => P(8)(74),s => s(8)(36),lamdaOut => P(7)(74));
G875: entity G port map(lamdaA => P(8)(73),lamdaB => P(8)(75),s => s(8)(37),lamdaOut => P(7)(75));
F876: entity F port map(lamdaA => P(8)(76),lamdaB => P(8)(78),lamdaOut => P(7)(76));
F877: entity F port map(lamdaA => P(8)(77),lamdaB => P(8)(79),lamdaOut => P(7)(77));
G878: entity G port map(lamdaA => P(8)(76),lamdaB => P(8)(78),s => s(8)(38),lamdaOut => P(7)(78));
G879: entity G port map(lamdaA => P(8)(77),lamdaB => P(8)(79),s => s(8)(39),lamdaOut => P(7)(79));
F880: entity F port map(lamdaA => P(8)(80),lamdaB => P(8)(82),lamdaOut => P(7)(80));
F881: entity F port map(lamdaA => P(8)(81),lamdaB => P(8)(83),lamdaOut => P(7)(81));
G882: entity G port map(lamdaA => P(8)(80),lamdaB => P(8)(82),s => s(8)(40),lamdaOut => P(7)(82));
G883: entity G port map(lamdaA => P(8)(81),lamdaB => P(8)(83),s => s(8)(41),lamdaOut => P(7)(83));
F884: entity F port map(lamdaA => P(8)(84),lamdaB => P(8)(86),lamdaOut => P(7)(84));
F885: entity F port map(lamdaA => P(8)(85),lamdaB => P(8)(87),lamdaOut => P(7)(85));
G886: entity G port map(lamdaA => P(8)(84),lamdaB => P(8)(86),s => s(8)(42),lamdaOut => P(7)(86));
G887: entity G port map(lamdaA => P(8)(85),lamdaB => P(8)(87),s => s(8)(43),lamdaOut => P(7)(87));
F888: entity F port map(lamdaA => P(8)(88),lamdaB => P(8)(90),lamdaOut => P(7)(88));
F889: entity F port map(lamdaA => P(8)(89),lamdaB => P(8)(91),lamdaOut => P(7)(89));
G890: entity G port map(lamdaA => P(8)(88),lamdaB => P(8)(90),s => s(8)(44),lamdaOut => P(7)(90));
G891: entity G port map(lamdaA => P(8)(89),lamdaB => P(8)(91),s => s(8)(45),lamdaOut => P(7)(91));
F892: entity F port map(lamdaA => P(8)(92),lamdaB => P(8)(94),lamdaOut => P(7)(92));
F893: entity F port map(lamdaA => P(8)(93),lamdaB => P(8)(95),lamdaOut => P(7)(93));
G894: entity G port map(lamdaA => P(8)(92),lamdaB => P(8)(94),s => s(8)(46),lamdaOut => P(7)(94));
G895: entity G port map(lamdaA => P(8)(93),lamdaB => P(8)(95),s => s(8)(47),lamdaOut => P(7)(95));
F896: entity F port map(lamdaA => P(8)(96),lamdaB => P(8)(98),lamdaOut => P(7)(96));
F897: entity F port map(lamdaA => P(8)(97),lamdaB => P(8)(99),lamdaOut => P(7)(97));
G898: entity G port map(lamdaA => P(8)(96),lamdaB => P(8)(98),s => s(8)(48),lamdaOut => P(7)(98));
G899: entity G port map(lamdaA => P(8)(97),lamdaB => P(8)(99),s => s(8)(49),lamdaOut => P(7)(99));
F8100: entity F port map(lamdaA => P(8)(100),lamdaB => P(8)(102),lamdaOut => P(7)(100));
F8101: entity F port map(lamdaA => P(8)(101),lamdaB => P(8)(103),lamdaOut => P(7)(101));
G8102: entity G port map(lamdaA => P(8)(100),lamdaB => P(8)(102),s => s(8)(50),lamdaOut => P(7)(102));
G8103: entity G port map(lamdaA => P(8)(101),lamdaB => P(8)(103),s => s(8)(51),lamdaOut => P(7)(103));
F8104: entity F port map(lamdaA => P(8)(104),lamdaB => P(8)(106),lamdaOut => P(7)(104));
F8105: entity F port map(lamdaA => P(8)(105),lamdaB => P(8)(107),lamdaOut => P(7)(105));
G8106: entity G port map(lamdaA => P(8)(104),lamdaB => P(8)(106),s => s(8)(52),lamdaOut => P(7)(106));
G8107: entity G port map(lamdaA => P(8)(105),lamdaB => P(8)(107),s => s(8)(53),lamdaOut => P(7)(107));
F8108: entity F port map(lamdaA => P(8)(108),lamdaB => P(8)(110),lamdaOut => P(7)(108));
F8109: entity F port map(lamdaA => P(8)(109),lamdaB => P(8)(111),lamdaOut => P(7)(109));
G8110: entity G port map(lamdaA => P(8)(108),lamdaB => P(8)(110),s => s(8)(54),lamdaOut => P(7)(110));
G8111: entity G port map(lamdaA => P(8)(109),lamdaB => P(8)(111),s => s(8)(55),lamdaOut => P(7)(111));
F8112: entity F port map(lamdaA => P(8)(112),lamdaB => P(8)(114),lamdaOut => P(7)(112));
F8113: entity F port map(lamdaA => P(8)(113),lamdaB => P(8)(115),lamdaOut => P(7)(113));
G8114: entity G port map(lamdaA => P(8)(112),lamdaB => P(8)(114),s => s(8)(56),lamdaOut => P(7)(114));
G8115: entity G port map(lamdaA => P(8)(113),lamdaB => P(8)(115),s => s(8)(57),lamdaOut => P(7)(115));
F8116: entity F port map(lamdaA => P(8)(116),lamdaB => P(8)(118),lamdaOut => P(7)(116));
F8117: entity F port map(lamdaA => P(8)(117),lamdaB => P(8)(119),lamdaOut => P(7)(117));
G8118: entity G port map(lamdaA => P(8)(116),lamdaB => P(8)(118),s => s(8)(58),lamdaOut => P(7)(118));
G8119: entity G port map(lamdaA => P(8)(117),lamdaB => P(8)(119),s => s(8)(59),lamdaOut => P(7)(119));
F8120: entity F port map(lamdaA => P(8)(120),lamdaB => P(8)(122),lamdaOut => P(7)(120));
F8121: entity F port map(lamdaA => P(8)(121),lamdaB => P(8)(123),lamdaOut => P(7)(121));
G8122: entity G port map(lamdaA => P(8)(120),lamdaB => P(8)(122),s => s(8)(60),lamdaOut => P(7)(122));
G8123: entity G port map(lamdaA => P(8)(121),lamdaB => P(8)(123),s => s(8)(61),lamdaOut => P(7)(123));
F8124: entity F port map(lamdaA => P(8)(124),lamdaB => P(8)(126),lamdaOut => P(7)(124));
F8125: entity F port map(lamdaA => P(8)(125),lamdaB => P(8)(127),lamdaOut => P(7)(125));
G8126: entity G port map(lamdaA => P(8)(124),lamdaB => P(8)(126),s => s(8)(62),lamdaOut => P(7)(126));
G8127: entity G port map(lamdaA => P(8)(125),lamdaB => P(8)(127),s => s(8)(63),lamdaOut => P(7)(127));
F8128: entity F port map(lamdaA => P(8)(128),lamdaB => P(8)(130),lamdaOut => P(7)(128));
F8129: entity F port map(lamdaA => P(8)(129),lamdaB => P(8)(131),lamdaOut => P(7)(129));
G8130: entity G port map(lamdaA => P(8)(128),lamdaB => P(8)(130),s => s(8)(64),lamdaOut => P(7)(130));
G8131: entity G port map(lamdaA => P(8)(129),lamdaB => P(8)(131),s => s(8)(65),lamdaOut => P(7)(131));
F8132: entity F port map(lamdaA => P(8)(132),lamdaB => P(8)(134),lamdaOut => P(7)(132));
F8133: entity F port map(lamdaA => P(8)(133),lamdaB => P(8)(135),lamdaOut => P(7)(133));
G8134: entity G port map(lamdaA => P(8)(132),lamdaB => P(8)(134),s => s(8)(66),lamdaOut => P(7)(134));
G8135: entity G port map(lamdaA => P(8)(133),lamdaB => P(8)(135),s => s(8)(67),lamdaOut => P(7)(135));
F8136: entity F port map(lamdaA => P(8)(136),lamdaB => P(8)(138),lamdaOut => P(7)(136));
F8137: entity F port map(lamdaA => P(8)(137),lamdaB => P(8)(139),lamdaOut => P(7)(137));
G8138: entity G port map(lamdaA => P(8)(136),lamdaB => P(8)(138),s => s(8)(68),lamdaOut => P(7)(138));
G8139: entity G port map(lamdaA => P(8)(137),lamdaB => P(8)(139),s => s(8)(69),lamdaOut => P(7)(139));
F8140: entity F port map(lamdaA => P(8)(140),lamdaB => P(8)(142),lamdaOut => P(7)(140));
F8141: entity F port map(lamdaA => P(8)(141),lamdaB => P(8)(143),lamdaOut => P(7)(141));
G8142: entity G port map(lamdaA => P(8)(140),lamdaB => P(8)(142),s => s(8)(70),lamdaOut => P(7)(142));
G8143: entity G port map(lamdaA => P(8)(141),lamdaB => P(8)(143),s => s(8)(71),lamdaOut => P(7)(143));
F8144: entity F port map(lamdaA => P(8)(144),lamdaB => P(8)(146),lamdaOut => P(7)(144));
F8145: entity F port map(lamdaA => P(8)(145),lamdaB => P(8)(147),lamdaOut => P(7)(145));
G8146: entity G port map(lamdaA => P(8)(144),lamdaB => P(8)(146),s => s(8)(72),lamdaOut => P(7)(146));
G8147: entity G port map(lamdaA => P(8)(145),lamdaB => P(8)(147),s => s(8)(73),lamdaOut => P(7)(147));
F8148: entity F port map(lamdaA => P(8)(148),lamdaB => P(8)(150),lamdaOut => P(7)(148));
F8149: entity F port map(lamdaA => P(8)(149),lamdaB => P(8)(151),lamdaOut => P(7)(149));
G8150: entity G port map(lamdaA => P(8)(148),lamdaB => P(8)(150),s => s(8)(74),lamdaOut => P(7)(150));
G8151: entity G port map(lamdaA => P(8)(149),lamdaB => P(8)(151),s => s(8)(75),lamdaOut => P(7)(151));
F8152: entity F port map(lamdaA => P(8)(152),lamdaB => P(8)(154),lamdaOut => P(7)(152));
F8153: entity F port map(lamdaA => P(8)(153),lamdaB => P(8)(155),lamdaOut => P(7)(153));
G8154: entity G port map(lamdaA => P(8)(152),lamdaB => P(8)(154),s => s(8)(76),lamdaOut => P(7)(154));
G8155: entity G port map(lamdaA => P(8)(153),lamdaB => P(8)(155),s => s(8)(77),lamdaOut => P(7)(155));
F8156: entity F port map(lamdaA => P(8)(156),lamdaB => P(8)(158),lamdaOut => P(7)(156));
F8157: entity F port map(lamdaA => P(8)(157),lamdaB => P(8)(159),lamdaOut => P(7)(157));
G8158: entity G port map(lamdaA => P(8)(156),lamdaB => P(8)(158),s => s(8)(78),lamdaOut => P(7)(158));
G8159: entity G port map(lamdaA => P(8)(157),lamdaB => P(8)(159),s => s(8)(79),lamdaOut => P(7)(159));
F8160: entity F port map(lamdaA => P(8)(160),lamdaB => P(8)(162),lamdaOut => P(7)(160));
F8161: entity F port map(lamdaA => P(8)(161),lamdaB => P(8)(163),lamdaOut => P(7)(161));
G8162: entity G port map(lamdaA => P(8)(160),lamdaB => P(8)(162),s => s(8)(80),lamdaOut => P(7)(162));
G8163: entity G port map(lamdaA => P(8)(161),lamdaB => P(8)(163),s => s(8)(81),lamdaOut => P(7)(163));
F8164: entity F port map(lamdaA => P(8)(164),lamdaB => P(8)(166),lamdaOut => P(7)(164));
F8165: entity F port map(lamdaA => P(8)(165),lamdaB => P(8)(167),lamdaOut => P(7)(165));
G8166: entity G port map(lamdaA => P(8)(164),lamdaB => P(8)(166),s => s(8)(82),lamdaOut => P(7)(166));
G8167: entity G port map(lamdaA => P(8)(165),lamdaB => P(8)(167),s => s(8)(83),lamdaOut => P(7)(167));
F8168: entity F port map(lamdaA => P(8)(168),lamdaB => P(8)(170),lamdaOut => P(7)(168));
F8169: entity F port map(lamdaA => P(8)(169),lamdaB => P(8)(171),lamdaOut => P(7)(169));
G8170: entity G port map(lamdaA => P(8)(168),lamdaB => P(8)(170),s => s(8)(84),lamdaOut => P(7)(170));
G8171: entity G port map(lamdaA => P(8)(169),lamdaB => P(8)(171),s => s(8)(85),lamdaOut => P(7)(171));
F8172: entity F port map(lamdaA => P(8)(172),lamdaB => P(8)(174),lamdaOut => P(7)(172));
F8173: entity F port map(lamdaA => P(8)(173),lamdaB => P(8)(175),lamdaOut => P(7)(173));
G8174: entity G port map(lamdaA => P(8)(172),lamdaB => P(8)(174),s => s(8)(86),lamdaOut => P(7)(174));
G8175: entity G port map(lamdaA => P(8)(173),lamdaB => P(8)(175),s => s(8)(87),lamdaOut => P(7)(175));
F8176: entity F port map(lamdaA => P(8)(176),lamdaB => P(8)(178),lamdaOut => P(7)(176));
F8177: entity F port map(lamdaA => P(8)(177),lamdaB => P(8)(179),lamdaOut => P(7)(177));
G8178: entity G port map(lamdaA => P(8)(176),lamdaB => P(8)(178),s => s(8)(88),lamdaOut => P(7)(178));
G8179: entity G port map(lamdaA => P(8)(177),lamdaB => P(8)(179),s => s(8)(89),lamdaOut => P(7)(179));
F8180: entity F port map(lamdaA => P(8)(180),lamdaB => P(8)(182),lamdaOut => P(7)(180));
F8181: entity F port map(lamdaA => P(8)(181),lamdaB => P(8)(183),lamdaOut => P(7)(181));
G8182: entity G port map(lamdaA => P(8)(180),lamdaB => P(8)(182),s => s(8)(90),lamdaOut => P(7)(182));
G8183: entity G port map(lamdaA => P(8)(181),lamdaB => P(8)(183),s => s(8)(91),lamdaOut => P(7)(183));
F8184: entity F port map(lamdaA => P(8)(184),lamdaB => P(8)(186),lamdaOut => P(7)(184));
F8185: entity F port map(lamdaA => P(8)(185),lamdaB => P(8)(187),lamdaOut => P(7)(185));
G8186: entity G port map(lamdaA => P(8)(184),lamdaB => P(8)(186),s => s(8)(92),lamdaOut => P(7)(186));
G8187: entity G port map(lamdaA => P(8)(185),lamdaB => P(8)(187),s => s(8)(93),lamdaOut => P(7)(187));
F8188: entity F port map(lamdaA => P(8)(188),lamdaB => P(8)(190),lamdaOut => P(7)(188));
F8189: entity F port map(lamdaA => P(8)(189),lamdaB => P(8)(191),lamdaOut => P(7)(189));
G8190: entity G port map(lamdaA => P(8)(188),lamdaB => P(8)(190),s => s(8)(94),lamdaOut => P(7)(190));
G8191: entity G port map(lamdaA => P(8)(189),lamdaB => P(8)(191),s => s(8)(95),lamdaOut => P(7)(191));
F8192: entity F port map(lamdaA => P(8)(192),lamdaB => P(8)(194),lamdaOut => P(7)(192));
F8193: entity F port map(lamdaA => P(8)(193),lamdaB => P(8)(195),lamdaOut => P(7)(193));
G8194: entity G port map(lamdaA => P(8)(192),lamdaB => P(8)(194),s => s(8)(96),lamdaOut => P(7)(194));
G8195: entity G port map(lamdaA => P(8)(193),lamdaB => P(8)(195),s => s(8)(97),lamdaOut => P(7)(195));
F8196: entity F port map(lamdaA => P(8)(196),lamdaB => P(8)(198),lamdaOut => P(7)(196));
F8197: entity F port map(lamdaA => P(8)(197),lamdaB => P(8)(199),lamdaOut => P(7)(197));
G8198: entity G port map(lamdaA => P(8)(196),lamdaB => P(8)(198),s => s(8)(98),lamdaOut => P(7)(198));
G8199: entity G port map(lamdaA => P(8)(197),lamdaB => P(8)(199),s => s(8)(99),lamdaOut => P(7)(199));
F8200: entity F port map(lamdaA => P(8)(200),lamdaB => P(8)(202),lamdaOut => P(7)(200));
F8201: entity F port map(lamdaA => P(8)(201),lamdaB => P(8)(203),lamdaOut => P(7)(201));
G8202: entity G port map(lamdaA => P(8)(200),lamdaB => P(8)(202),s => s(8)(100),lamdaOut => P(7)(202));
G8203: entity G port map(lamdaA => P(8)(201),lamdaB => P(8)(203),s => s(8)(101),lamdaOut => P(7)(203));
F8204: entity F port map(lamdaA => P(8)(204),lamdaB => P(8)(206),lamdaOut => P(7)(204));
F8205: entity F port map(lamdaA => P(8)(205),lamdaB => P(8)(207),lamdaOut => P(7)(205));
G8206: entity G port map(lamdaA => P(8)(204),lamdaB => P(8)(206),s => s(8)(102),lamdaOut => P(7)(206));
G8207: entity G port map(lamdaA => P(8)(205),lamdaB => P(8)(207),s => s(8)(103),lamdaOut => P(7)(207));
F8208: entity F port map(lamdaA => P(8)(208),lamdaB => P(8)(210),lamdaOut => P(7)(208));
F8209: entity F port map(lamdaA => P(8)(209),lamdaB => P(8)(211),lamdaOut => P(7)(209));
G8210: entity G port map(lamdaA => P(8)(208),lamdaB => P(8)(210),s => s(8)(104),lamdaOut => P(7)(210));
G8211: entity G port map(lamdaA => P(8)(209),lamdaB => P(8)(211),s => s(8)(105),lamdaOut => P(7)(211));
F8212: entity F port map(lamdaA => P(8)(212),lamdaB => P(8)(214),lamdaOut => P(7)(212));
F8213: entity F port map(lamdaA => P(8)(213),lamdaB => P(8)(215),lamdaOut => P(7)(213));
G8214: entity G port map(lamdaA => P(8)(212),lamdaB => P(8)(214),s => s(8)(106),lamdaOut => P(7)(214));
G8215: entity G port map(lamdaA => P(8)(213),lamdaB => P(8)(215),s => s(8)(107),lamdaOut => P(7)(215));
F8216: entity F port map(lamdaA => P(8)(216),lamdaB => P(8)(218),lamdaOut => P(7)(216));
F8217: entity F port map(lamdaA => P(8)(217),lamdaB => P(8)(219),lamdaOut => P(7)(217));
G8218: entity G port map(lamdaA => P(8)(216),lamdaB => P(8)(218),s => s(8)(108),lamdaOut => P(7)(218));
G8219: entity G port map(lamdaA => P(8)(217),lamdaB => P(8)(219),s => s(8)(109),lamdaOut => P(7)(219));
F8220: entity F port map(lamdaA => P(8)(220),lamdaB => P(8)(222),lamdaOut => P(7)(220));
F8221: entity F port map(lamdaA => P(8)(221),lamdaB => P(8)(223),lamdaOut => P(7)(221));
G8222: entity G port map(lamdaA => P(8)(220),lamdaB => P(8)(222),s => s(8)(110),lamdaOut => P(7)(222));
G8223: entity G port map(lamdaA => P(8)(221),lamdaB => P(8)(223),s => s(8)(111),lamdaOut => P(7)(223));
F8224: entity F port map(lamdaA => P(8)(224),lamdaB => P(8)(226),lamdaOut => P(7)(224));
F8225: entity F port map(lamdaA => P(8)(225),lamdaB => P(8)(227),lamdaOut => P(7)(225));
G8226: entity G port map(lamdaA => P(8)(224),lamdaB => P(8)(226),s => s(8)(112),lamdaOut => P(7)(226));
G8227: entity G port map(lamdaA => P(8)(225),lamdaB => P(8)(227),s => s(8)(113),lamdaOut => P(7)(227));
F8228: entity F port map(lamdaA => P(8)(228),lamdaB => P(8)(230),lamdaOut => P(7)(228));
F8229: entity F port map(lamdaA => P(8)(229),lamdaB => P(8)(231),lamdaOut => P(7)(229));
G8230: entity G port map(lamdaA => P(8)(228),lamdaB => P(8)(230),s => s(8)(114),lamdaOut => P(7)(230));
G8231: entity G port map(lamdaA => P(8)(229),lamdaB => P(8)(231),s => s(8)(115),lamdaOut => P(7)(231));
F8232: entity F port map(lamdaA => P(8)(232),lamdaB => P(8)(234),lamdaOut => P(7)(232));
F8233: entity F port map(lamdaA => P(8)(233),lamdaB => P(8)(235),lamdaOut => P(7)(233));
G8234: entity G port map(lamdaA => P(8)(232),lamdaB => P(8)(234),s => s(8)(116),lamdaOut => P(7)(234));
G8235: entity G port map(lamdaA => P(8)(233),lamdaB => P(8)(235),s => s(8)(117),lamdaOut => P(7)(235));
F8236: entity F port map(lamdaA => P(8)(236),lamdaB => P(8)(238),lamdaOut => P(7)(236));
F8237: entity F port map(lamdaA => P(8)(237),lamdaB => P(8)(239),lamdaOut => P(7)(237));
G8238: entity G port map(lamdaA => P(8)(236),lamdaB => P(8)(238),s => s(8)(118),lamdaOut => P(7)(238));
G8239: entity G port map(lamdaA => P(8)(237),lamdaB => P(8)(239),s => s(8)(119),lamdaOut => P(7)(239));
F8240: entity F port map(lamdaA => P(8)(240),lamdaB => P(8)(242),lamdaOut => P(7)(240));
F8241: entity F port map(lamdaA => P(8)(241),lamdaB => P(8)(243),lamdaOut => P(7)(241));
G8242: entity G port map(lamdaA => P(8)(240),lamdaB => P(8)(242),s => s(8)(120),lamdaOut => P(7)(242));
G8243: entity G port map(lamdaA => P(8)(241),lamdaB => P(8)(243),s => s(8)(121),lamdaOut => P(7)(243));
F8244: entity F port map(lamdaA => P(8)(244),lamdaB => P(8)(246),lamdaOut => P(7)(244));
F8245: entity F port map(lamdaA => P(8)(245),lamdaB => P(8)(247),lamdaOut => P(7)(245));
G8246: entity G port map(lamdaA => P(8)(244),lamdaB => P(8)(246),s => s(8)(122),lamdaOut => P(7)(246));
G8247: entity G port map(lamdaA => P(8)(245),lamdaB => P(8)(247),s => s(8)(123),lamdaOut => P(7)(247));
F8248: entity F port map(lamdaA => P(8)(248),lamdaB => P(8)(250),lamdaOut => P(7)(248));
F8249: entity F port map(lamdaA => P(8)(249),lamdaB => P(8)(251),lamdaOut => P(7)(249));
G8250: entity G port map(lamdaA => P(8)(248),lamdaB => P(8)(250),s => s(8)(124),lamdaOut => P(7)(250));
G8251: entity G port map(lamdaA => P(8)(249),lamdaB => P(8)(251),s => s(8)(125),lamdaOut => P(7)(251));
F8252: entity F port map(lamdaA => P(8)(252),lamdaB => P(8)(254),lamdaOut => P(7)(252));
F8253: entity F port map(lamdaA => P(8)(253),lamdaB => P(8)(255),lamdaOut => P(7)(253));
G8254: entity G port map(lamdaA => P(8)(252),lamdaB => P(8)(254),s => s(8)(126),lamdaOut => P(7)(254));
G8255: entity G port map(lamdaA => P(8)(253),lamdaB => P(8)(255),s => s(8)(127),lamdaOut => P(7)(255));
F8256: entity F port map(lamdaA => P(8)(256),lamdaB => P(8)(258),lamdaOut => P(7)(256));
F8257: entity F port map(lamdaA => P(8)(257),lamdaB => P(8)(259),lamdaOut => P(7)(257));
G8258: entity G port map(lamdaA => P(8)(256),lamdaB => P(8)(258),s => s(8)(128),lamdaOut => P(7)(258));
G8259: entity G port map(lamdaA => P(8)(257),lamdaB => P(8)(259),s => s(8)(129),lamdaOut => P(7)(259));
F8260: entity F port map(lamdaA => P(8)(260),lamdaB => P(8)(262),lamdaOut => P(7)(260));
F8261: entity F port map(lamdaA => P(8)(261),lamdaB => P(8)(263),lamdaOut => P(7)(261));
G8262: entity G port map(lamdaA => P(8)(260),lamdaB => P(8)(262),s => s(8)(130),lamdaOut => P(7)(262));
G8263: entity G port map(lamdaA => P(8)(261),lamdaB => P(8)(263),s => s(8)(131),lamdaOut => P(7)(263));
F8264: entity F port map(lamdaA => P(8)(264),lamdaB => P(8)(266),lamdaOut => P(7)(264));
F8265: entity F port map(lamdaA => P(8)(265),lamdaB => P(8)(267),lamdaOut => P(7)(265));
G8266: entity G port map(lamdaA => P(8)(264),lamdaB => P(8)(266),s => s(8)(132),lamdaOut => P(7)(266));
G8267: entity G port map(lamdaA => P(8)(265),lamdaB => P(8)(267),s => s(8)(133),lamdaOut => P(7)(267));
F8268: entity F port map(lamdaA => P(8)(268),lamdaB => P(8)(270),lamdaOut => P(7)(268));
F8269: entity F port map(lamdaA => P(8)(269),lamdaB => P(8)(271),lamdaOut => P(7)(269));
G8270: entity G port map(lamdaA => P(8)(268),lamdaB => P(8)(270),s => s(8)(134),lamdaOut => P(7)(270));
G8271: entity G port map(lamdaA => P(8)(269),lamdaB => P(8)(271),s => s(8)(135),lamdaOut => P(7)(271));
F8272: entity F port map(lamdaA => P(8)(272),lamdaB => P(8)(274),lamdaOut => P(7)(272));
F8273: entity F port map(lamdaA => P(8)(273),lamdaB => P(8)(275),lamdaOut => P(7)(273));
G8274: entity G port map(lamdaA => P(8)(272),lamdaB => P(8)(274),s => s(8)(136),lamdaOut => P(7)(274));
G8275: entity G port map(lamdaA => P(8)(273),lamdaB => P(8)(275),s => s(8)(137),lamdaOut => P(7)(275));
F8276: entity F port map(lamdaA => P(8)(276),lamdaB => P(8)(278),lamdaOut => P(7)(276));
F8277: entity F port map(lamdaA => P(8)(277),lamdaB => P(8)(279),lamdaOut => P(7)(277));
G8278: entity G port map(lamdaA => P(8)(276),lamdaB => P(8)(278),s => s(8)(138),lamdaOut => P(7)(278));
G8279: entity G port map(lamdaA => P(8)(277),lamdaB => P(8)(279),s => s(8)(139),lamdaOut => P(7)(279));
F8280: entity F port map(lamdaA => P(8)(280),lamdaB => P(8)(282),lamdaOut => P(7)(280));
F8281: entity F port map(lamdaA => P(8)(281),lamdaB => P(8)(283),lamdaOut => P(7)(281));
G8282: entity G port map(lamdaA => P(8)(280),lamdaB => P(8)(282),s => s(8)(140),lamdaOut => P(7)(282));
G8283: entity G port map(lamdaA => P(8)(281),lamdaB => P(8)(283),s => s(8)(141),lamdaOut => P(7)(283));
F8284: entity F port map(lamdaA => P(8)(284),lamdaB => P(8)(286),lamdaOut => P(7)(284));
F8285: entity F port map(lamdaA => P(8)(285),lamdaB => P(8)(287),lamdaOut => P(7)(285));
G8286: entity G port map(lamdaA => P(8)(284),lamdaB => P(8)(286),s => s(8)(142),lamdaOut => P(7)(286));
G8287: entity G port map(lamdaA => P(8)(285),lamdaB => P(8)(287),s => s(8)(143),lamdaOut => P(7)(287));
F8288: entity F port map(lamdaA => P(8)(288),lamdaB => P(8)(290),lamdaOut => P(7)(288));
F8289: entity F port map(lamdaA => P(8)(289),lamdaB => P(8)(291),lamdaOut => P(7)(289));
G8290: entity G port map(lamdaA => P(8)(288),lamdaB => P(8)(290),s => s(8)(144),lamdaOut => P(7)(290));
G8291: entity G port map(lamdaA => P(8)(289),lamdaB => P(8)(291),s => s(8)(145),lamdaOut => P(7)(291));
F8292: entity F port map(lamdaA => P(8)(292),lamdaB => P(8)(294),lamdaOut => P(7)(292));
F8293: entity F port map(lamdaA => P(8)(293),lamdaB => P(8)(295),lamdaOut => P(7)(293));
G8294: entity G port map(lamdaA => P(8)(292),lamdaB => P(8)(294),s => s(8)(146),lamdaOut => P(7)(294));
G8295: entity G port map(lamdaA => P(8)(293),lamdaB => P(8)(295),s => s(8)(147),lamdaOut => P(7)(295));
F8296: entity F port map(lamdaA => P(8)(296),lamdaB => P(8)(298),lamdaOut => P(7)(296));
F8297: entity F port map(lamdaA => P(8)(297),lamdaB => P(8)(299),lamdaOut => P(7)(297));
G8298: entity G port map(lamdaA => P(8)(296),lamdaB => P(8)(298),s => s(8)(148),lamdaOut => P(7)(298));
G8299: entity G port map(lamdaA => P(8)(297),lamdaB => P(8)(299),s => s(8)(149),lamdaOut => P(7)(299));
F8300: entity F port map(lamdaA => P(8)(300),lamdaB => P(8)(302),lamdaOut => P(7)(300));
F8301: entity F port map(lamdaA => P(8)(301),lamdaB => P(8)(303),lamdaOut => P(7)(301));
G8302: entity G port map(lamdaA => P(8)(300),lamdaB => P(8)(302),s => s(8)(150),lamdaOut => P(7)(302));
G8303: entity G port map(lamdaA => P(8)(301),lamdaB => P(8)(303),s => s(8)(151),lamdaOut => P(7)(303));
F8304: entity F port map(lamdaA => P(8)(304),lamdaB => P(8)(306),lamdaOut => P(7)(304));
F8305: entity F port map(lamdaA => P(8)(305),lamdaB => P(8)(307),lamdaOut => P(7)(305));
G8306: entity G port map(lamdaA => P(8)(304),lamdaB => P(8)(306),s => s(8)(152),lamdaOut => P(7)(306));
G8307: entity G port map(lamdaA => P(8)(305),lamdaB => P(8)(307),s => s(8)(153),lamdaOut => P(7)(307));
F8308: entity F port map(lamdaA => P(8)(308),lamdaB => P(8)(310),lamdaOut => P(7)(308));
F8309: entity F port map(lamdaA => P(8)(309),lamdaB => P(8)(311),lamdaOut => P(7)(309));
G8310: entity G port map(lamdaA => P(8)(308),lamdaB => P(8)(310),s => s(8)(154),lamdaOut => P(7)(310));
G8311: entity G port map(lamdaA => P(8)(309),lamdaB => P(8)(311),s => s(8)(155),lamdaOut => P(7)(311));
F8312: entity F port map(lamdaA => P(8)(312),lamdaB => P(8)(314),lamdaOut => P(7)(312));
F8313: entity F port map(lamdaA => P(8)(313),lamdaB => P(8)(315),lamdaOut => P(7)(313));
G8314: entity G port map(lamdaA => P(8)(312),lamdaB => P(8)(314),s => s(8)(156),lamdaOut => P(7)(314));
G8315: entity G port map(lamdaA => P(8)(313),lamdaB => P(8)(315),s => s(8)(157),lamdaOut => P(7)(315));
F8316: entity F port map(lamdaA => P(8)(316),lamdaB => P(8)(318),lamdaOut => P(7)(316));
F8317: entity F port map(lamdaA => P(8)(317),lamdaB => P(8)(319),lamdaOut => P(7)(317));
G8318: entity G port map(lamdaA => P(8)(316),lamdaB => P(8)(318),s => s(8)(158),lamdaOut => P(7)(318));
G8319: entity G port map(lamdaA => P(8)(317),lamdaB => P(8)(319),s => s(8)(159),lamdaOut => P(7)(319));
F8320: entity F port map(lamdaA => P(8)(320),lamdaB => P(8)(322),lamdaOut => P(7)(320));
F8321: entity F port map(lamdaA => P(8)(321),lamdaB => P(8)(323),lamdaOut => P(7)(321));
G8322: entity G port map(lamdaA => P(8)(320),lamdaB => P(8)(322),s => s(8)(160),lamdaOut => P(7)(322));
G8323: entity G port map(lamdaA => P(8)(321),lamdaB => P(8)(323),s => s(8)(161),lamdaOut => P(7)(323));
F8324: entity F port map(lamdaA => P(8)(324),lamdaB => P(8)(326),lamdaOut => P(7)(324));
F8325: entity F port map(lamdaA => P(8)(325),lamdaB => P(8)(327),lamdaOut => P(7)(325));
G8326: entity G port map(lamdaA => P(8)(324),lamdaB => P(8)(326),s => s(8)(162),lamdaOut => P(7)(326));
G8327: entity G port map(lamdaA => P(8)(325),lamdaB => P(8)(327),s => s(8)(163),lamdaOut => P(7)(327));
F8328: entity F port map(lamdaA => P(8)(328),lamdaB => P(8)(330),lamdaOut => P(7)(328));
F8329: entity F port map(lamdaA => P(8)(329),lamdaB => P(8)(331),lamdaOut => P(7)(329));
G8330: entity G port map(lamdaA => P(8)(328),lamdaB => P(8)(330),s => s(8)(164),lamdaOut => P(7)(330));
G8331: entity G port map(lamdaA => P(8)(329),lamdaB => P(8)(331),s => s(8)(165),lamdaOut => P(7)(331));
F8332: entity F port map(lamdaA => P(8)(332),lamdaB => P(8)(334),lamdaOut => P(7)(332));
F8333: entity F port map(lamdaA => P(8)(333),lamdaB => P(8)(335),lamdaOut => P(7)(333));
G8334: entity G port map(lamdaA => P(8)(332),lamdaB => P(8)(334),s => s(8)(166),lamdaOut => P(7)(334));
G8335: entity G port map(lamdaA => P(8)(333),lamdaB => P(8)(335),s => s(8)(167),lamdaOut => P(7)(335));
F8336: entity F port map(lamdaA => P(8)(336),lamdaB => P(8)(338),lamdaOut => P(7)(336));
F8337: entity F port map(lamdaA => P(8)(337),lamdaB => P(8)(339),lamdaOut => P(7)(337));
G8338: entity G port map(lamdaA => P(8)(336),lamdaB => P(8)(338),s => s(8)(168),lamdaOut => P(7)(338));
G8339: entity G port map(lamdaA => P(8)(337),lamdaB => P(8)(339),s => s(8)(169),lamdaOut => P(7)(339));
F8340: entity F port map(lamdaA => P(8)(340),lamdaB => P(8)(342),lamdaOut => P(7)(340));
F8341: entity F port map(lamdaA => P(8)(341),lamdaB => P(8)(343),lamdaOut => P(7)(341));
G8342: entity G port map(lamdaA => P(8)(340),lamdaB => P(8)(342),s => s(8)(170),lamdaOut => P(7)(342));
G8343: entity G port map(lamdaA => P(8)(341),lamdaB => P(8)(343),s => s(8)(171),lamdaOut => P(7)(343));
F8344: entity F port map(lamdaA => P(8)(344),lamdaB => P(8)(346),lamdaOut => P(7)(344));
F8345: entity F port map(lamdaA => P(8)(345),lamdaB => P(8)(347),lamdaOut => P(7)(345));
G8346: entity G port map(lamdaA => P(8)(344),lamdaB => P(8)(346),s => s(8)(172),lamdaOut => P(7)(346));
G8347: entity G port map(lamdaA => P(8)(345),lamdaB => P(8)(347),s => s(8)(173),lamdaOut => P(7)(347));
F8348: entity F port map(lamdaA => P(8)(348),lamdaB => P(8)(350),lamdaOut => P(7)(348));
F8349: entity F port map(lamdaA => P(8)(349),lamdaB => P(8)(351),lamdaOut => P(7)(349));
G8350: entity G port map(lamdaA => P(8)(348),lamdaB => P(8)(350),s => s(8)(174),lamdaOut => P(7)(350));
G8351: entity G port map(lamdaA => P(8)(349),lamdaB => P(8)(351),s => s(8)(175),lamdaOut => P(7)(351));
F8352: entity F port map(lamdaA => P(8)(352),lamdaB => P(8)(354),lamdaOut => P(7)(352));
F8353: entity F port map(lamdaA => P(8)(353),lamdaB => P(8)(355),lamdaOut => P(7)(353));
G8354: entity G port map(lamdaA => P(8)(352),lamdaB => P(8)(354),s => s(8)(176),lamdaOut => P(7)(354));
G8355: entity G port map(lamdaA => P(8)(353),lamdaB => P(8)(355),s => s(8)(177),lamdaOut => P(7)(355));
F8356: entity F port map(lamdaA => P(8)(356),lamdaB => P(8)(358),lamdaOut => P(7)(356));
F8357: entity F port map(lamdaA => P(8)(357),lamdaB => P(8)(359),lamdaOut => P(7)(357));
G8358: entity G port map(lamdaA => P(8)(356),lamdaB => P(8)(358),s => s(8)(178),lamdaOut => P(7)(358));
G8359: entity G port map(lamdaA => P(8)(357),lamdaB => P(8)(359),s => s(8)(179),lamdaOut => P(7)(359));
F8360: entity F port map(lamdaA => P(8)(360),lamdaB => P(8)(362),lamdaOut => P(7)(360));
F8361: entity F port map(lamdaA => P(8)(361),lamdaB => P(8)(363),lamdaOut => P(7)(361));
G8362: entity G port map(lamdaA => P(8)(360),lamdaB => P(8)(362),s => s(8)(180),lamdaOut => P(7)(362));
G8363: entity G port map(lamdaA => P(8)(361),lamdaB => P(8)(363),s => s(8)(181),lamdaOut => P(7)(363));
F8364: entity F port map(lamdaA => P(8)(364),lamdaB => P(8)(366),lamdaOut => P(7)(364));
F8365: entity F port map(lamdaA => P(8)(365),lamdaB => P(8)(367),lamdaOut => P(7)(365));
G8366: entity G port map(lamdaA => P(8)(364),lamdaB => P(8)(366),s => s(8)(182),lamdaOut => P(7)(366));
G8367: entity G port map(lamdaA => P(8)(365),lamdaB => P(8)(367),s => s(8)(183),lamdaOut => P(7)(367));
F8368: entity F port map(lamdaA => P(8)(368),lamdaB => P(8)(370),lamdaOut => P(7)(368));
F8369: entity F port map(lamdaA => P(8)(369),lamdaB => P(8)(371),lamdaOut => P(7)(369));
G8370: entity G port map(lamdaA => P(8)(368),lamdaB => P(8)(370),s => s(8)(184),lamdaOut => P(7)(370));
G8371: entity G port map(lamdaA => P(8)(369),lamdaB => P(8)(371),s => s(8)(185),lamdaOut => P(7)(371));
F8372: entity F port map(lamdaA => P(8)(372),lamdaB => P(8)(374),lamdaOut => P(7)(372));
F8373: entity F port map(lamdaA => P(8)(373),lamdaB => P(8)(375),lamdaOut => P(7)(373));
G8374: entity G port map(lamdaA => P(8)(372),lamdaB => P(8)(374),s => s(8)(186),lamdaOut => P(7)(374));
G8375: entity G port map(lamdaA => P(8)(373),lamdaB => P(8)(375),s => s(8)(187),lamdaOut => P(7)(375));
F8376: entity F port map(lamdaA => P(8)(376),lamdaB => P(8)(378),lamdaOut => P(7)(376));
F8377: entity F port map(lamdaA => P(8)(377),lamdaB => P(8)(379),lamdaOut => P(7)(377));
G8378: entity G port map(lamdaA => P(8)(376),lamdaB => P(8)(378),s => s(8)(188),lamdaOut => P(7)(378));
G8379: entity G port map(lamdaA => P(8)(377),lamdaB => P(8)(379),s => s(8)(189),lamdaOut => P(7)(379));
F8380: entity F port map(lamdaA => P(8)(380),lamdaB => P(8)(382),lamdaOut => P(7)(380));
F8381: entity F port map(lamdaA => P(8)(381),lamdaB => P(8)(383),lamdaOut => P(7)(381));
G8382: entity G port map(lamdaA => P(8)(380),lamdaB => P(8)(382),s => s(8)(190),lamdaOut => P(7)(382));
G8383: entity G port map(lamdaA => P(8)(381),lamdaB => P(8)(383),s => s(8)(191),lamdaOut => P(7)(383));
F8384: entity F port map(lamdaA => P(8)(384),lamdaB => P(8)(386),lamdaOut => P(7)(384));
F8385: entity F port map(lamdaA => P(8)(385),lamdaB => P(8)(387),lamdaOut => P(7)(385));
G8386: entity G port map(lamdaA => P(8)(384),lamdaB => P(8)(386),s => s(8)(192),lamdaOut => P(7)(386));
G8387: entity G port map(lamdaA => P(8)(385),lamdaB => P(8)(387),s => s(8)(193),lamdaOut => P(7)(387));
F8388: entity F port map(lamdaA => P(8)(388),lamdaB => P(8)(390),lamdaOut => P(7)(388));
F8389: entity F port map(lamdaA => P(8)(389),lamdaB => P(8)(391),lamdaOut => P(7)(389));
G8390: entity G port map(lamdaA => P(8)(388),lamdaB => P(8)(390),s => s(8)(194),lamdaOut => P(7)(390));
G8391: entity G port map(lamdaA => P(8)(389),lamdaB => P(8)(391),s => s(8)(195),lamdaOut => P(7)(391));
F8392: entity F port map(lamdaA => P(8)(392),lamdaB => P(8)(394),lamdaOut => P(7)(392));
F8393: entity F port map(lamdaA => P(8)(393),lamdaB => P(8)(395),lamdaOut => P(7)(393));
G8394: entity G port map(lamdaA => P(8)(392),lamdaB => P(8)(394),s => s(8)(196),lamdaOut => P(7)(394));
G8395: entity G port map(lamdaA => P(8)(393),lamdaB => P(8)(395),s => s(8)(197),lamdaOut => P(7)(395));
F8396: entity F port map(lamdaA => P(8)(396),lamdaB => P(8)(398),lamdaOut => P(7)(396));
F8397: entity F port map(lamdaA => P(8)(397),lamdaB => P(8)(399),lamdaOut => P(7)(397));
G8398: entity G port map(lamdaA => P(8)(396),lamdaB => P(8)(398),s => s(8)(198),lamdaOut => P(7)(398));
G8399: entity G port map(lamdaA => P(8)(397),lamdaB => P(8)(399),s => s(8)(199),lamdaOut => P(7)(399));
F8400: entity F port map(lamdaA => P(8)(400),lamdaB => P(8)(402),lamdaOut => P(7)(400));
F8401: entity F port map(lamdaA => P(8)(401),lamdaB => P(8)(403),lamdaOut => P(7)(401));
G8402: entity G port map(lamdaA => P(8)(400),lamdaB => P(8)(402),s => s(8)(200),lamdaOut => P(7)(402));
G8403: entity G port map(lamdaA => P(8)(401),lamdaB => P(8)(403),s => s(8)(201),lamdaOut => P(7)(403));
F8404: entity F port map(lamdaA => P(8)(404),lamdaB => P(8)(406),lamdaOut => P(7)(404));
F8405: entity F port map(lamdaA => P(8)(405),lamdaB => P(8)(407),lamdaOut => P(7)(405));
G8406: entity G port map(lamdaA => P(8)(404),lamdaB => P(8)(406),s => s(8)(202),lamdaOut => P(7)(406));
G8407: entity G port map(lamdaA => P(8)(405),lamdaB => P(8)(407),s => s(8)(203),lamdaOut => P(7)(407));
F8408: entity F port map(lamdaA => P(8)(408),lamdaB => P(8)(410),lamdaOut => P(7)(408));
F8409: entity F port map(lamdaA => P(8)(409),lamdaB => P(8)(411),lamdaOut => P(7)(409));
G8410: entity G port map(lamdaA => P(8)(408),lamdaB => P(8)(410),s => s(8)(204),lamdaOut => P(7)(410));
G8411: entity G port map(lamdaA => P(8)(409),lamdaB => P(8)(411),s => s(8)(205),lamdaOut => P(7)(411));
F8412: entity F port map(lamdaA => P(8)(412),lamdaB => P(8)(414),lamdaOut => P(7)(412));
F8413: entity F port map(lamdaA => P(8)(413),lamdaB => P(8)(415),lamdaOut => P(7)(413));
G8414: entity G port map(lamdaA => P(8)(412),lamdaB => P(8)(414),s => s(8)(206),lamdaOut => P(7)(414));
G8415: entity G port map(lamdaA => P(8)(413),lamdaB => P(8)(415),s => s(8)(207),lamdaOut => P(7)(415));
F8416: entity F port map(lamdaA => P(8)(416),lamdaB => P(8)(418),lamdaOut => P(7)(416));
F8417: entity F port map(lamdaA => P(8)(417),lamdaB => P(8)(419),lamdaOut => P(7)(417));
G8418: entity G port map(lamdaA => P(8)(416),lamdaB => P(8)(418),s => s(8)(208),lamdaOut => P(7)(418));
G8419: entity G port map(lamdaA => P(8)(417),lamdaB => P(8)(419),s => s(8)(209),lamdaOut => P(7)(419));
F8420: entity F port map(lamdaA => P(8)(420),lamdaB => P(8)(422),lamdaOut => P(7)(420));
F8421: entity F port map(lamdaA => P(8)(421),lamdaB => P(8)(423),lamdaOut => P(7)(421));
G8422: entity G port map(lamdaA => P(8)(420),lamdaB => P(8)(422),s => s(8)(210),lamdaOut => P(7)(422));
G8423: entity G port map(lamdaA => P(8)(421),lamdaB => P(8)(423),s => s(8)(211),lamdaOut => P(7)(423));
F8424: entity F port map(lamdaA => P(8)(424),lamdaB => P(8)(426),lamdaOut => P(7)(424));
F8425: entity F port map(lamdaA => P(8)(425),lamdaB => P(8)(427),lamdaOut => P(7)(425));
G8426: entity G port map(lamdaA => P(8)(424),lamdaB => P(8)(426),s => s(8)(212),lamdaOut => P(7)(426));
G8427: entity G port map(lamdaA => P(8)(425),lamdaB => P(8)(427),s => s(8)(213),lamdaOut => P(7)(427));
F8428: entity F port map(lamdaA => P(8)(428),lamdaB => P(8)(430),lamdaOut => P(7)(428));
F8429: entity F port map(lamdaA => P(8)(429),lamdaB => P(8)(431),lamdaOut => P(7)(429));
G8430: entity G port map(lamdaA => P(8)(428),lamdaB => P(8)(430),s => s(8)(214),lamdaOut => P(7)(430));
G8431: entity G port map(lamdaA => P(8)(429),lamdaB => P(8)(431),s => s(8)(215),lamdaOut => P(7)(431));
F8432: entity F port map(lamdaA => P(8)(432),lamdaB => P(8)(434),lamdaOut => P(7)(432));
F8433: entity F port map(lamdaA => P(8)(433),lamdaB => P(8)(435),lamdaOut => P(7)(433));
G8434: entity G port map(lamdaA => P(8)(432),lamdaB => P(8)(434),s => s(8)(216),lamdaOut => P(7)(434));
G8435: entity G port map(lamdaA => P(8)(433),lamdaB => P(8)(435),s => s(8)(217),lamdaOut => P(7)(435));
F8436: entity F port map(lamdaA => P(8)(436),lamdaB => P(8)(438),lamdaOut => P(7)(436));
F8437: entity F port map(lamdaA => P(8)(437),lamdaB => P(8)(439),lamdaOut => P(7)(437));
G8438: entity G port map(lamdaA => P(8)(436),lamdaB => P(8)(438),s => s(8)(218),lamdaOut => P(7)(438));
G8439: entity G port map(lamdaA => P(8)(437),lamdaB => P(8)(439),s => s(8)(219),lamdaOut => P(7)(439));
F8440: entity F port map(lamdaA => P(8)(440),lamdaB => P(8)(442),lamdaOut => P(7)(440));
F8441: entity F port map(lamdaA => P(8)(441),lamdaB => P(8)(443),lamdaOut => P(7)(441));
G8442: entity G port map(lamdaA => P(8)(440),lamdaB => P(8)(442),s => s(8)(220),lamdaOut => P(7)(442));
G8443: entity G port map(lamdaA => P(8)(441),lamdaB => P(8)(443),s => s(8)(221),lamdaOut => P(7)(443));
F8444: entity F port map(lamdaA => P(8)(444),lamdaB => P(8)(446),lamdaOut => P(7)(444));
F8445: entity F port map(lamdaA => P(8)(445),lamdaB => P(8)(447),lamdaOut => P(7)(445));
G8446: entity G port map(lamdaA => P(8)(444),lamdaB => P(8)(446),s => s(8)(222),lamdaOut => P(7)(446));
G8447: entity G port map(lamdaA => P(8)(445),lamdaB => P(8)(447),s => s(8)(223),lamdaOut => P(7)(447));
F8448: entity F port map(lamdaA => P(8)(448),lamdaB => P(8)(450),lamdaOut => P(7)(448));
F8449: entity F port map(lamdaA => P(8)(449),lamdaB => P(8)(451),lamdaOut => P(7)(449));
G8450: entity G port map(lamdaA => P(8)(448),lamdaB => P(8)(450),s => s(8)(224),lamdaOut => P(7)(450));
G8451: entity G port map(lamdaA => P(8)(449),lamdaB => P(8)(451),s => s(8)(225),lamdaOut => P(7)(451));
F8452: entity F port map(lamdaA => P(8)(452),lamdaB => P(8)(454),lamdaOut => P(7)(452));
F8453: entity F port map(lamdaA => P(8)(453),lamdaB => P(8)(455),lamdaOut => P(7)(453));
G8454: entity G port map(lamdaA => P(8)(452),lamdaB => P(8)(454),s => s(8)(226),lamdaOut => P(7)(454));
G8455: entity G port map(lamdaA => P(8)(453),lamdaB => P(8)(455),s => s(8)(227),lamdaOut => P(7)(455));
F8456: entity F port map(lamdaA => P(8)(456),lamdaB => P(8)(458),lamdaOut => P(7)(456));
F8457: entity F port map(lamdaA => P(8)(457),lamdaB => P(8)(459),lamdaOut => P(7)(457));
G8458: entity G port map(lamdaA => P(8)(456),lamdaB => P(8)(458),s => s(8)(228),lamdaOut => P(7)(458));
G8459: entity G port map(lamdaA => P(8)(457),lamdaB => P(8)(459),s => s(8)(229),lamdaOut => P(7)(459));
F8460: entity F port map(lamdaA => P(8)(460),lamdaB => P(8)(462),lamdaOut => P(7)(460));
F8461: entity F port map(lamdaA => P(8)(461),lamdaB => P(8)(463),lamdaOut => P(7)(461));
G8462: entity G port map(lamdaA => P(8)(460),lamdaB => P(8)(462),s => s(8)(230),lamdaOut => P(7)(462));
G8463: entity G port map(lamdaA => P(8)(461),lamdaB => P(8)(463),s => s(8)(231),lamdaOut => P(7)(463));
F8464: entity F port map(lamdaA => P(8)(464),lamdaB => P(8)(466),lamdaOut => P(7)(464));
F8465: entity F port map(lamdaA => P(8)(465),lamdaB => P(8)(467),lamdaOut => P(7)(465));
G8466: entity G port map(lamdaA => P(8)(464),lamdaB => P(8)(466),s => s(8)(232),lamdaOut => P(7)(466));
G8467: entity G port map(lamdaA => P(8)(465),lamdaB => P(8)(467),s => s(8)(233),lamdaOut => P(7)(467));
F8468: entity F port map(lamdaA => P(8)(468),lamdaB => P(8)(470),lamdaOut => P(7)(468));
F8469: entity F port map(lamdaA => P(8)(469),lamdaB => P(8)(471),lamdaOut => P(7)(469));
G8470: entity G port map(lamdaA => P(8)(468),lamdaB => P(8)(470),s => s(8)(234),lamdaOut => P(7)(470));
G8471: entity G port map(lamdaA => P(8)(469),lamdaB => P(8)(471),s => s(8)(235),lamdaOut => P(7)(471));
F8472: entity F port map(lamdaA => P(8)(472),lamdaB => P(8)(474),lamdaOut => P(7)(472));
F8473: entity F port map(lamdaA => P(8)(473),lamdaB => P(8)(475),lamdaOut => P(7)(473));
G8474: entity G port map(lamdaA => P(8)(472),lamdaB => P(8)(474),s => s(8)(236),lamdaOut => P(7)(474));
G8475: entity G port map(lamdaA => P(8)(473),lamdaB => P(8)(475),s => s(8)(237),lamdaOut => P(7)(475));
F8476: entity F port map(lamdaA => P(8)(476),lamdaB => P(8)(478),lamdaOut => P(7)(476));
F8477: entity F port map(lamdaA => P(8)(477),lamdaB => P(8)(479),lamdaOut => P(7)(477));
G8478: entity G port map(lamdaA => P(8)(476),lamdaB => P(8)(478),s => s(8)(238),lamdaOut => P(7)(478));
G8479: entity G port map(lamdaA => P(8)(477),lamdaB => P(8)(479),s => s(8)(239),lamdaOut => P(7)(479));
F8480: entity F port map(lamdaA => P(8)(480),lamdaB => P(8)(482),lamdaOut => P(7)(480));
F8481: entity F port map(lamdaA => P(8)(481),lamdaB => P(8)(483),lamdaOut => P(7)(481));
G8482: entity G port map(lamdaA => P(8)(480),lamdaB => P(8)(482),s => s(8)(240),lamdaOut => P(7)(482));
G8483: entity G port map(lamdaA => P(8)(481),lamdaB => P(8)(483),s => s(8)(241),lamdaOut => P(7)(483));
F8484: entity F port map(lamdaA => P(8)(484),lamdaB => P(8)(486),lamdaOut => P(7)(484));
F8485: entity F port map(lamdaA => P(8)(485),lamdaB => P(8)(487),lamdaOut => P(7)(485));
G8486: entity G port map(lamdaA => P(8)(484),lamdaB => P(8)(486),s => s(8)(242),lamdaOut => P(7)(486));
G8487: entity G port map(lamdaA => P(8)(485),lamdaB => P(8)(487),s => s(8)(243),lamdaOut => P(7)(487));
F8488: entity F port map(lamdaA => P(8)(488),lamdaB => P(8)(490),lamdaOut => P(7)(488));
F8489: entity F port map(lamdaA => P(8)(489),lamdaB => P(8)(491),lamdaOut => P(7)(489));
G8490: entity G port map(lamdaA => P(8)(488),lamdaB => P(8)(490),s => s(8)(244),lamdaOut => P(7)(490));
G8491: entity G port map(lamdaA => P(8)(489),lamdaB => P(8)(491),s => s(8)(245),lamdaOut => P(7)(491));
F8492: entity F port map(lamdaA => P(8)(492),lamdaB => P(8)(494),lamdaOut => P(7)(492));
F8493: entity F port map(lamdaA => P(8)(493),lamdaB => P(8)(495),lamdaOut => P(7)(493));
G8494: entity G port map(lamdaA => P(8)(492),lamdaB => P(8)(494),s => s(8)(246),lamdaOut => P(7)(494));
G8495: entity G port map(lamdaA => P(8)(493),lamdaB => P(8)(495),s => s(8)(247),lamdaOut => P(7)(495));
F8496: entity F port map(lamdaA => P(8)(496),lamdaB => P(8)(498),lamdaOut => P(7)(496));
F8497: entity F port map(lamdaA => P(8)(497),lamdaB => P(8)(499),lamdaOut => P(7)(497));
G8498: entity G port map(lamdaA => P(8)(496),lamdaB => P(8)(498),s => s(8)(248),lamdaOut => P(7)(498));
G8499: entity G port map(lamdaA => P(8)(497),lamdaB => P(8)(499),s => s(8)(249),lamdaOut => P(7)(499));
F8500: entity F port map(lamdaA => P(8)(500),lamdaB => P(8)(502),lamdaOut => P(7)(500));
F8501: entity F port map(lamdaA => P(8)(501),lamdaB => P(8)(503),lamdaOut => P(7)(501));
G8502: entity G port map(lamdaA => P(8)(500),lamdaB => P(8)(502),s => s(8)(250),lamdaOut => P(7)(502));
G8503: entity G port map(lamdaA => P(8)(501),lamdaB => P(8)(503),s => s(8)(251),lamdaOut => P(7)(503));
F8504: entity F port map(lamdaA => P(8)(504),lamdaB => P(8)(506),lamdaOut => P(7)(504));
F8505: entity F port map(lamdaA => P(8)(505),lamdaB => P(8)(507),lamdaOut => P(7)(505));
G8506: entity G port map(lamdaA => P(8)(504),lamdaB => P(8)(506),s => s(8)(252),lamdaOut => P(7)(506));
G8507: entity G port map(lamdaA => P(8)(505),lamdaB => P(8)(507),s => s(8)(253),lamdaOut => P(7)(507));
F8508: entity F port map(lamdaA => P(8)(508),lamdaB => P(8)(510),lamdaOut => P(7)(508));
F8509: entity F port map(lamdaA => P(8)(509),lamdaB => P(8)(511),lamdaOut => P(7)(509));
G8510: entity G port map(lamdaA => P(8)(508),lamdaB => P(8)(510),s => s(8)(254),lamdaOut => P(7)(510));
G8511: entity G port map(lamdaA => P(8)(509),lamdaB => P(8)(511),s => s(8)(255),lamdaOut => P(7)(511));
-- STAGE 7
F70: entity F port map(lamdaA => P(7)(0),lamdaB => P(7)(4),lamdaOut => P(6)(0));
F71: entity F port map(lamdaA => P(7)(1),lamdaB => P(7)(5),lamdaOut => P(6)(1));
F72: entity F port map(lamdaA => P(7)(2),lamdaB => P(7)(6),lamdaOut => P(6)(2));
F73: entity F port map(lamdaA => P(7)(3),lamdaB => P(7)(7),lamdaOut => P(6)(3));
G74: entity G port map(lamdaA => P(7)(0),lamdaB => P(7)(4),s => s(7)(0),lamdaOut => P(6)(4));
G75: entity G port map(lamdaA => P(7)(1),lamdaB => P(7)(5),s => s(7)(1),lamdaOut => P(6)(5));
G76: entity G port map(lamdaA => P(7)(2),lamdaB => P(7)(6),s => s(7)(2),lamdaOut => P(6)(6));
G77: entity G port map(lamdaA => P(7)(3),lamdaB => P(7)(7),s => s(7)(3),lamdaOut => P(6)(7));
F78: entity F port map(lamdaA => P(7)(8),lamdaB => P(7)(12),lamdaOut => P(6)(8));
F79: entity F port map(lamdaA => P(7)(9),lamdaB => P(7)(13),lamdaOut => P(6)(9));
F710: entity F port map(lamdaA => P(7)(10),lamdaB => P(7)(14),lamdaOut => P(6)(10));
F711: entity F port map(lamdaA => P(7)(11),lamdaB => P(7)(15),lamdaOut => P(6)(11));
G712: entity G port map(lamdaA => P(7)(8),lamdaB => P(7)(12),s => s(7)(4),lamdaOut => P(6)(12));
G713: entity G port map(lamdaA => P(7)(9),lamdaB => P(7)(13),s => s(7)(5),lamdaOut => P(6)(13));
G714: entity G port map(lamdaA => P(7)(10),lamdaB => P(7)(14),s => s(7)(6),lamdaOut => P(6)(14));
G715: entity G port map(lamdaA => P(7)(11),lamdaB => P(7)(15),s => s(7)(7),lamdaOut => P(6)(15));
F716: entity F port map(lamdaA => P(7)(16),lamdaB => P(7)(20),lamdaOut => P(6)(16));
F717: entity F port map(lamdaA => P(7)(17),lamdaB => P(7)(21),lamdaOut => P(6)(17));
F718: entity F port map(lamdaA => P(7)(18),lamdaB => P(7)(22),lamdaOut => P(6)(18));
F719: entity F port map(lamdaA => P(7)(19),lamdaB => P(7)(23),lamdaOut => P(6)(19));
G720: entity G port map(lamdaA => P(7)(16),lamdaB => P(7)(20),s => s(7)(8),lamdaOut => P(6)(20));
G721: entity G port map(lamdaA => P(7)(17),lamdaB => P(7)(21),s => s(7)(9),lamdaOut => P(6)(21));
G722: entity G port map(lamdaA => P(7)(18),lamdaB => P(7)(22),s => s(7)(10),lamdaOut => P(6)(22));
G723: entity G port map(lamdaA => P(7)(19),lamdaB => P(7)(23),s => s(7)(11),lamdaOut => P(6)(23));
F724: entity F port map(lamdaA => P(7)(24),lamdaB => P(7)(28),lamdaOut => P(6)(24));
F725: entity F port map(lamdaA => P(7)(25),lamdaB => P(7)(29),lamdaOut => P(6)(25));
F726: entity F port map(lamdaA => P(7)(26),lamdaB => P(7)(30),lamdaOut => P(6)(26));
F727: entity F port map(lamdaA => P(7)(27),lamdaB => P(7)(31),lamdaOut => P(6)(27));
G728: entity G port map(lamdaA => P(7)(24),lamdaB => P(7)(28),s => s(7)(12),lamdaOut => P(6)(28));
G729: entity G port map(lamdaA => P(7)(25),lamdaB => P(7)(29),s => s(7)(13),lamdaOut => P(6)(29));
G730: entity G port map(lamdaA => P(7)(26),lamdaB => P(7)(30),s => s(7)(14),lamdaOut => P(6)(30));
G731: entity G port map(lamdaA => P(7)(27),lamdaB => P(7)(31),s => s(7)(15),lamdaOut => P(6)(31));
F732: entity F port map(lamdaA => P(7)(32),lamdaB => P(7)(36),lamdaOut => P(6)(32));
F733: entity F port map(lamdaA => P(7)(33),lamdaB => P(7)(37),lamdaOut => P(6)(33));
F734: entity F port map(lamdaA => P(7)(34),lamdaB => P(7)(38),lamdaOut => P(6)(34));
F735: entity F port map(lamdaA => P(7)(35),lamdaB => P(7)(39),lamdaOut => P(6)(35));
G736: entity G port map(lamdaA => P(7)(32),lamdaB => P(7)(36),s => s(7)(16),lamdaOut => P(6)(36));
G737: entity G port map(lamdaA => P(7)(33),lamdaB => P(7)(37),s => s(7)(17),lamdaOut => P(6)(37));
G738: entity G port map(lamdaA => P(7)(34),lamdaB => P(7)(38),s => s(7)(18),lamdaOut => P(6)(38));
G739: entity G port map(lamdaA => P(7)(35),lamdaB => P(7)(39),s => s(7)(19),lamdaOut => P(6)(39));
F740: entity F port map(lamdaA => P(7)(40),lamdaB => P(7)(44),lamdaOut => P(6)(40));
F741: entity F port map(lamdaA => P(7)(41),lamdaB => P(7)(45),lamdaOut => P(6)(41));
F742: entity F port map(lamdaA => P(7)(42),lamdaB => P(7)(46),lamdaOut => P(6)(42));
F743: entity F port map(lamdaA => P(7)(43),lamdaB => P(7)(47),lamdaOut => P(6)(43));
G744: entity G port map(lamdaA => P(7)(40),lamdaB => P(7)(44),s => s(7)(20),lamdaOut => P(6)(44));
G745: entity G port map(lamdaA => P(7)(41),lamdaB => P(7)(45),s => s(7)(21),lamdaOut => P(6)(45));
G746: entity G port map(lamdaA => P(7)(42),lamdaB => P(7)(46),s => s(7)(22),lamdaOut => P(6)(46));
G747: entity G port map(lamdaA => P(7)(43),lamdaB => P(7)(47),s => s(7)(23),lamdaOut => P(6)(47));
F748: entity F port map(lamdaA => P(7)(48),lamdaB => P(7)(52),lamdaOut => P(6)(48));
F749: entity F port map(lamdaA => P(7)(49),lamdaB => P(7)(53),lamdaOut => P(6)(49));
F750: entity F port map(lamdaA => P(7)(50),lamdaB => P(7)(54),lamdaOut => P(6)(50));
F751: entity F port map(lamdaA => P(7)(51),lamdaB => P(7)(55),lamdaOut => P(6)(51));
G752: entity G port map(lamdaA => P(7)(48),lamdaB => P(7)(52),s => s(7)(24),lamdaOut => P(6)(52));
G753: entity G port map(lamdaA => P(7)(49),lamdaB => P(7)(53),s => s(7)(25),lamdaOut => P(6)(53));
G754: entity G port map(lamdaA => P(7)(50),lamdaB => P(7)(54),s => s(7)(26),lamdaOut => P(6)(54));
G755: entity G port map(lamdaA => P(7)(51),lamdaB => P(7)(55),s => s(7)(27),lamdaOut => P(6)(55));
F756: entity F port map(lamdaA => P(7)(56),lamdaB => P(7)(60),lamdaOut => P(6)(56));
F757: entity F port map(lamdaA => P(7)(57),lamdaB => P(7)(61),lamdaOut => P(6)(57));
F758: entity F port map(lamdaA => P(7)(58),lamdaB => P(7)(62),lamdaOut => P(6)(58));
F759: entity F port map(lamdaA => P(7)(59),lamdaB => P(7)(63),lamdaOut => P(6)(59));
G760: entity G port map(lamdaA => P(7)(56),lamdaB => P(7)(60),s => s(7)(28),lamdaOut => P(6)(60));
G761: entity G port map(lamdaA => P(7)(57),lamdaB => P(7)(61),s => s(7)(29),lamdaOut => P(6)(61));
G762: entity G port map(lamdaA => P(7)(58),lamdaB => P(7)(62),s => s(7)(30),lamdaOut => P(6)(62));
G763: entity G port map(lamdaA => P(7)(59),lamdaB => P(7)(63),s => s(7)(31),lamdaOut => P(6)(63));
F764: entity F port map(lamdaA => P(7)(64),lamdaB => P(7)(68),lamdaOut => P(6)(64));
F765: entity F port map(lamdaA => P(7)(65),lamdaB => P(7)(69),lamdaOut => P(6)(65));
F766: entity F port map(lamdaA => P(7)(66),lamdaB => P(7)(70),lamdaOut => P(6)(66));
F767: entity F port map(lamdaA => P(7)(67),lamdaB => P(7)(71),lamdaOut => P(6)(67));
G768: entity G port map(lamdaA => P(7)(64),lamdaB => P(7)(68),s => s(7)(32),lamdaOut => P(6)(68));
G769: entity G port map(lamdaA => P(7)(65),lamdaB => P(7)(69),s => s(7)(33),lamdaOut => P(6)(69));
G770: entity G port map(lamdaA => P(7)(66),lamdaB => P(7)(70),s => s(7)(34),lamdaOut => P(6)(70));
G771: entity G port map(lamdaA => P(7)(67),lamdaB => P(7)(71),s => s(7)(35),lamdaOut => P(6)(71));
F772: entity F port map(lamdaA => P(7)(72),lamdaB => P(7)(76),lamdaOut => P(6)(72));
F773: entity F port map(lamdaA => P(7)(73),lamdaB => P(7)(77),lamdaOut => P(6)(73));
F774: entity F port map(lamdaA => P(7)(74),lamdaB => P(7)(78),lamdaOut => P(6)(74));
F775: entity F port map(lamdaA => P(7)(75),lamdaB => P(7)(79),lamdaOut => P(6)(75));
G776: entity G port map(lamdaA => P(7)(72),lamdaB => P(7)(76),s => s(7)(36),lamdaOut => P(6)(76));
G777: entity G port map(lamdaA => P(7)(73),lamdaB => P(7)(77),s => s(7)(37),lamdaOut => P(6)(77));
G778: entity G port map(lamdaA => P(7)(74),lamdaB => P(7)(78),s => s(7)(38),lamdaOut => P(6)(78));
G779: entity G port map(lamdaA => P(7)(75),lamdaB => P(7)(79),s => s(7)(39),lamdaOut => P(6)(79));
F780: entity F port map(lamdaA => P(7)(80),lamdaB => P(7)(84),lamdaOut => P(6)(80));
F781: entity F port map(lamdaA => P(7)(81),lamdaB => P(7)(85),lamdaOut => P(6)(81));
F782: entity F port map(lamdaA => P(7)(82),lamdaB => P(7)(86),lamdaOut => P(6)(82));
F783: entity F port map(lamdaA => P(7)(83),lamdaB => P(7)(87),lamdaOut => P(6)(83));
G784: entity G port map(lamdaA => P(7)(80),lamdaB => P(7)(84),s => s(7)(40),lamdaOut => P(6)(84));
G785: entity G port map(lamdaA => P(7)(81),lamdaB => P(7)(85),s => s(7)(41),lamdaOut => P(6)(85));
G786: entity G port map(lamdaA => P(7)(82),lamdaB => P(7)(86),s => s(7)(42),lamdaOut => P(6)(86));
G787: entity G port map(lamdaA => P(7)(83),lamdaB => P(7)(87),s => s(7)(43),lamdaOut => P(6)(87));
F788: entity F port map(lamdaA => P(7)(88),lamdaB => P(7)(92),lamdaOut => P(6)(88));
F789: entity F port map(lamdaA => P(7)(89),lamdaB => P(7)(93),lamdaOut => P(6)(89));
F790: entity F port map(lamdaA => P(7)(90),lamdaB => P(7)(94),lamdaOut => P(6)(90));
F791: entity F port map(lamdaA => P(7)(91),lamdaB => P(7)(95),lamdaOut => P(6)(91));
G792: entity G port map(lamdaA => P(7)(88),lamdaB => P(7)(92),s => s(7)(44),lamdaOut => P(6)(92));
G793: entity G port map(lamdaA => P(7)(89),lamdaB => P(7)(93),s => s(7)(45),lamdaOut => P(6)(93));
G794: entity G port map(lamdaA => P(7)(90),lamdaB => P(7)(94),s => s(7)(46),lamdaOut => P(6)(94));
G795: entity G port map(lamdaA => P(7)(91),lamdaB => P(7)(95),s => s(7)(47),lamdaOut => P(6)(95));
F796: entity F port map(lamdaA => P(7)(96),lamdaB => P(7)(100),lamdaOut => P(6)(96));
F797: entity F port map(lamdaA => P(7)(97),lamdaB => P(7)(101),lamdaOut => P(6)(97));
F798: entity F port map(lamdaA => P(7)(98),lamdaB => P(7)(102),lamdaOut => P(6)(98));
F799: entity F port map(lamdaA => P(7)(99),lamdaB => P(7)(103),lamdaOut => P(6)(99));
G7100: entity G port map(lamdaA => P(7)(96),lamdaB => P(7)(100),s => s(7)(48),lamdaOut => P(6)(100));
G7101: entity G port map(lamdaA => P(7)(97),lamdaB => P(7)(101),s => s(7)(49),lamdaOut => P(6)(101));
G7102: entity G port map(lamdaA => P(7)(98),lamdaB => P(7)(102),s => s(7)(50),lamdaOut => P(6)(102));
G7103: entity G port map(lamdaA => P(7)(99),lamdaB => P(7)(103),s => s(7)(51),lamdaOut => P(6)(103));
F7104: entity F port map(lamdaA => P(7)(104),lamdaB => P(7)(108),lamdaOut => P(6)(104));
F7105: entity F port map(lamdaA => P(7)(105),lamdaB => P(7)(109),lamdaOut => P(6)(105));
F7106: entity F port map(lamdaA => P(7)(106),lamdaB => P(7)(110),lamdaOut => P(6)(106));
F7107: entity F port map(lamdaA => P(7)(107),lamdaB => P(7)(111),lamdaOut => P(6)(107));
G7108: entity G port map(lamdaA => P(7)(104),lamdaB => P(7)(108),s => s(7)(52),lamdaOut => P(6)(108));
G7109: entity G port map(lamdaA => P(7)(105),lamdaB => P(7)(109),s => s(7)(53),lamdaOut => P(6)(109));
G7110: entity G port map(lamdaA => P(7)(106),lamdaB => P(7)(110),s => s(7)(54),lamdaOut => P(6)(110));
G7111: entity G port map(lamdaA => P(7)(107),lamdaB => P(7)(111),s => s(7)(55),lamdaOut => P(6)(111));
F7112: entity F port map(lamdaA => P(7)(112),lamdaB => P(7)(116),lamdaOut => P(6)(112));
F7113: entity F port map(lamdaA => P(7)(113),lamdaB => P(7)(117),lamdaOut => P(6)(113));
F7114: entity F port map(lamdaA => P(7)(114),lamdaB => P(7)(118),lamdaOut => P(6)(114));
F7115: entity F port map(lamdaA => P(7)(115),lamdaB => P(7)(119),lamdaOut => P(6)(115));
G7116: entity G port map(lamdaA => P(7)(112),lamdaB => P(7)(116),s => s(7)(56),lamdaOut => P(6)(116));
G7117: entity G port map(lamdaA => P(7)(113),lamdaB => P(7)(117),s => s(7)(57),lamdaOut => P(6)(117));
G7118: entity G port map(lamdaA => P(7)(114),lamdaB => P(7)(118),s => s(7)(58),lamdaOut => P(6)(118));
G7119: entity G port map(lamdaA => P(7)(115),lamdaB => P(7)(119),s => s(7)(59),lamdaOut => P(6)(119));
F7120: entity F port map(lamdaA => P(7)(120),lamdaB => P(7)(124),lamdaOut => P(6)(120));
F7121: entity F port map(lamdaA => P(7)(121),lamdaB => P(7)(125),lamdaOut => P(6)(121));
F7122: entity F port map(lamdaA => P(7)(122),lamdaB => P(7)(126),lamdaOut => P(6)(122));
F7123: entity F port map(lamdaA => P(7)(123),lamdaB => P(7)(127),lamdaOut => P(6)(123));
G7124: entity G port map(lamdaA => P(7)(120),lamdaB => P(7)(124),s => s(7)(60),lamdaOut => P(6)(124));
G7125: entity G port map(lamdaA => P(7)(121),lamdaB => P(7)(125),s => s(7)(61),lamdaOut => P(6)(125));
G7126: entity G port map(lamdaA => P(7)(122),lamdaB => P(7)(126),s => s(7)(62),lamdaOut => P(6)(126));
G7127: entity G port map(lamdaA => P(7)(123),lamdaB => P(7)(127),s => s(7)(63),lamdaOut => P(6)(127));
F7128: entity F port map(lamdaA => P(7)(128),lamdaB => P(7)(132),lamdaOut => P(6)(128));
F7129: entity F port map(lamdaA => P(7)(129),lamdaB => P(7)(133),lamdaOut => P(6)(129));
F7130: entity F port map(lamdaA => P(7)(130),lamdaB => P(7)(134),lamdaOut => P(6)(130));
F7131: entity F port map(lamdaA => P(7)(131),lamdaB => P(7)(135),lamdaOut => P(6)(131));
G7132: entity G port map(lamdaA => P(7)(128),lamdaB => P(7)(132),s => s(7)(64),lamdaOut => P(6)(132));
G7133: entity G port map(lamdaA => P(7)(129),lamdaB => P(7)(133),s => s(7)(65),lamdaOut => P(6)(133));
G7134: entity G port map(lamdaA => P(7)(130),lamdaB => P(7)(134),s => s(7)(66),lamdaOut => P(6)(134));
G7135: entity G port map(lamdaA => P(7)(131),lamdaB => P(7)(135),s => s(7)(67),lamdaOut => P(6)(135));
F7136: entity F port map(lamdaA => P(7)(136),lamdaB => P(7)(140),lamdaOut => P(6)(136));
F7137: entity F port map(lamdaA => P(7)(137),lamdaB => P(7)(141),lamdaOut => P(6)(137));
F7138: entity F port map(lamdaA => P(7)(138),lamdaB => P(7)(142),lamdaOut => P(6)(138));
F7139: entity F port map(lamdaA => P(7)(139),lamdaB => P(7)(143),lamdaOut => P(6)(139));
G7140: entity G port map(lamdaA => P(7)(136),lamdaB => P(7)(140),s => s(7)(68),lamdaOut => P(6)(140));
G7141: entity G port map(lamdaA => P(7)(137),lamdaB => P(7)(141),s => s(7)(69),lamdaOut => P(6)(141));
G7142: entity G port map(lamdaA => P(7)(138),lamdaB => P(7)(142),s => s(7)(70),lamdaOut => P(6)(142));
G7143: entity G port map(lamdaA => P(7)(139),lamdaB => P(7)(143),s => s(7)(71),lamdaOut => P(6)(143));
F7144: entity F port map(lamdaA => P(7)(144),lamdaB => P(7)(148),lamdaOut => P(6)(144));
F7145: entity F port map(lamdaA => P(7)(145),lamdaB => P(7)(149),lamdaOut => P(6)(145));
F7146: entity F port map(lamdaA => P(7)(146),lamdaB => P(7)(150),lamdaOut => P(6)(146));
F7147: entity F port map(lamdaA => P(7)(147),lamdaB => P(7)(151),lamdaOut => P(6)(147));
G7148: entity G port map(lamdaA => P(7)(144),lamdaB => P(7)(148),s => s(7)(72),lamdaOut => P(6)(148));
G7149: entity G port map(lamdaA => P(7)(145),lamdaB => P(7)(149),s => s(7)(73),lamdaOut => P(6)(149));
G7150: entity G port map(lamdaA => P(7)(146),lamdaB => P(7)(150),s => s(7)(74),lamdaOut => P(6)(150));
G7151: entity G port map(lamdaA => P(7)(147),lamdaB => P(7)(151),s => s(7)(75),lamdaOut => P(6)(151));
F7152: entity F port map(lamdaA => P(7)(152),lamdaB => P(7)(156),lamdaOut => P(6)(152));
F7153: entity F port map(lamdaA => P(7)(153),lamdaB => P(7)(157),lamdaOut => P(6)(153));
F7154: entity F port map(lamdaA => P(7)(154),lamdaB => P(7)(158),lamdaOut => P(6)(154));
F7155: entity F port map(lamdaA => P(7)(155),lamdaB => P(7)(159),lamdaOut => P(6)(155));
G7156: entity G port map(lamdaA => P(7)(152),lamdaB => P(7)(156),s => s(7)(76),lamdaOut => P(6)(156));
G7157: entity G port map(lamdaA => P(7)(153),lamdaB => P(7)(157),s => s(7)(77),lamdaOut => P(6)(157));
G7158: entity G port map(lamdaA => P(7)(154),lamdaB => P(7)(158),s => s(7)(78),lamdaOut => P(6)(158));
G7159: entity G port map(lamdaA => P(7)(155),lamdaB => P(7)(159),s => s(7)(79),lamdaOut => P(6)(159));
F7160: entity F port map(lamdaA => P(7)(160),lamdaB => P(7)(164),lamdaOut => P(6)(160));
F7161: entity F port map(lamdaA => P(7)(161),lamdaB => P(7)(165),lamdaOut => P(6)(161));
F7162: entity F port map(lamdaA => P(7)(162),lamdaB => P(7)(166),lamdaOut => P(6)(162));
F7163: entity F port map(lamdaA => P(7)(163),lamdaB => P(7)(167),lamdaOut => P(6)(163));
G7164: entity G port map(lamdaA => P(7)(160),lamdaB => P(7)(164),s => s(7)(80),lamdaOut => P(6)(164));
G7165: entity G port map(lamdaA => P(7)(161),lamdaB => P(7)(165),s => s(7)(81),lamdaOut => P(6)(165));
G7166: entity G port map(lamdaA => P(7)(162),lamdaB => P(7)(166),s => s(7)(82),lamdaOut => P(6)(166));
G7167: entity G port map(lamdaA => P(7)(163),lamdaB => P(7)(167),s => s(7)(83),lamdaOut => P(6)(167));
F7168: entity F port map(lamdaA => P(7)(168),lamdaB => P(7)(172),lamdaOut => P(6)(168));
F7169: entity F port map(lamdaA => P(7)(169),lamdaB => P(7)(173),lamdaOut => P(6)(169));
F7170: entity F port map(lamdaA => P(7)(170),lamdaB => P(7)(174),lamdaOut => P(6)(170));
F7171: entity F port map(lamdaA => P(7)(171),lamdaB => P(7)(175),lamdaOut => P(6)(171));
G7172: entity G port map(lamdaA => P(7)(168),lamdaB => P(7)(172),s => s(7)(84),lamdaOut => P(6)(172));
G7173: entity G port map(lamdaA => P(7)(169),lamdaB => P(7)(173),s => s(7)(85),lamdaOut => P(6)(173));
G7174: entity G port map(lamdaA => P(7)(170),lamdaB => P(7)(174),s => s(7)(86),lamdaOut => P(6)(174));
G7175: entity G port map(lamdaA => P(7)(171),lamdaB => P(7)(175),s => s(7)(87),lamdaOut => P(6)(175));
F7176: entity F port map(lamdaA => P(7)(176),lamdaB => P(7)(180),lamdaOut => P(6)(176));
F7177: entity F port map(lamdaA => P(7)(177),lamdaB => P(7)(181),lamdaOut => P(6)(177));
F7178: entity F port map(lamdaA => P(7)(178),lamdaB => P(7)(182),lamdaOut => P(6)(178));
F7179: entity F port map(lamdaA => P(7)(179),lamdaB => P(7)(183),lamdaOut => P(6)(179));
G7180: entity G port map(lamdaA => P(7)(176),lamdaB => P(7)(180),s => s(7)(88),lamdaOut => P(6)(180));
G7181: entity G port map(lamdaA => P(7)(177),lamdaB => P(7)(181),s => s(7)(89),lamdaOut => P(6)(181));
G7182: entity G port map(lamdaA => P(7)(178),lamdaB => P(7)(182),s => s(7)(90),lamdaOut => P(6)(182));
G7183: entity G port map(lamdaA => P(7)(179),lamdaB => P(7)(183),s => s(7)(91),lamdaOut => P(6)(183));
F7184: entity F port map(lamdaA => P(7)(184),lamdaB => P(7)(188),lamdaOut => P(6)(184));
F7185: entity F port map(lamdaA => P(7)(185),lamdaB => P(7)(189),lamdaOut => P(6)(185));
F7186: entity F port map(lamdaA => P(7)(186),lamdaB => P(7)(190),lamdaOut => P(6)(186));
F7187: entity F port map(lamdaA => P(7)(187),lamdaB => P(7)(191),lamdaOut => P(6)(187));
G7188: entity G port map(lamdaA => P(7)(184),lamdaB => P(7)(188),s => s(7)(92),lamdaOut => P(6)(188));
G7189: entity G port map(lamdaA => P(7)(185),lamdaB => P(7)(189),s => s(7)(93),lamdaOut => P(6)(189));
G7190: entity G port map(lamdaA => P(7)(186),lamdaB => P(7)(190),s => s(7)(94),lamdaOut => P(6)(190));
G7191: entity G port map(lamdaA => P(7)(187),lamdaB => P(7)(191),s => s(7)(95),lamdaOut => P(6)(191));
F7192: entity F port map(lamdaA => P(7)(192),lamdaB => P(7)(196),lamdaOut => P(6)(192));
F7193: entity F port map(lamdaA => P(7)(193),lamdaB => P(7)(197),lamdaOut => P(6)(193));
F7194: entity F port map(lamdaA => P(7)(194),lamdaB => P(7)(198),lamdaOut => P(6)(194));
F7195: entity F port map(lamdaA => P(7)(195),lamdaB => P(7)(199),lamdaOut => P(6)(195));
G7196: entity G port map(lamdaA => P(7)(192),lamdaB => P(7)(196),s => s(7)(96),lamdaOut => P(6)(196));
G7197: entity G port map(lamdaA => P(7)(193),lamdaB => P(7)(197),s => s(7)(97),lamdaOut => P(6)(197));
G7198: entity G port map(lamdaA => P(7)(194),lamdaB => P(7)(198),s => s(7)(98),lamdaOut => P(6)(198));
G7199: entity G port map(lamdaA => P(7)(195),lamdaB => P(7)(199),s => s(7)(99),lamdaOut => P(6)(199));
F7200: entity F port map(lamdaA => P(7)(200),lamdaB => P(7)(204),lamdaOut => P(6)(200));
F7201: entity F port map(lamdaA => P(7)(201),lamdaB => P(7)(205),lamdaOut => P(6)(201));
F7202: entity F port map(lamdaA => P(7)(202),lamdaB => P(7)(206),lamdaOut => P(6)(202));
F7203: entity F port map(lamdaA => P(7)(203),lamdaB => P(7)(207),lamdaOut => P(6)(203));
G7204: entity G port map(lamdaA => P(7)(200),lamdaB => P(7)(204),s => s(7)(100),lamdaOut => P(6)(204));
G7205: entity G port map(lamdaA => P(7)(201),lamdaB => P(7)(205),s => s(7)(101),lamdaOut => P(6)(205));
G7206: entity G port map(lamdaA => P(7)(202),lamdaB => P(7)(206),s => s(7)(102),lamdaOut => P(6)(206));
G7207: entity G port map(lamdaA => P(7)(203),lamdaB => P(7)(207),s => s(7)(103),lamdaOut => P(6)(207));
F7208: entity F port map(lamdaA => P(7)(208),lamdaB => P(7)(212),lamdaOut => P(6)(208));
F7209: entity F port map(lamdaA => P(7)(209),lamdaB => P(7)(213),lamdaOut => P(6)(209));
F7210: entity F port map(lamdaA => P(7)(210),lamdaB => P(7)(214),lamdaOut => P(6)(210));
F7211: entity F port map(lamdaA => P(7)(211),lamdaB => P(7)(215),lamdaOut => P(6)(211));
G7212: entity G port map(lamdaA => P(7)(208),lamdaB => P(7)(212),s => s(7)(104),lamdaOut => P(6)(212));
G7213: entity G port map(lamdaA => P(7)(209),lamdaB => P(7)(213),s => s(7)(105),lamdaOut => P(6)(213));
G7214: entity G port map(lamdaA => P(7)(210),lamdaB => P(7)(214),s => s(7)(106),lamdaOut => P(6)(214));
G7215: entity G port map(lamdaA => P(7)(211),lamdaB => P(7)(215),s => s(7)(107),lamdaOut => P(6)(215));
F7216: entity F port map(lamdaA => P(7)(216),lamdaB => P(7)(220),lamdaOut => P(6)(216));
F7217: entity F port map(lamdaA => P(7)(217),lamdaB => P(7)(221),lamdaOut => P(6)(217));
F7218: entity F port map(lamdaA => P(7)(218),lamdaB => P(7)(222),lamdaOut => P(6)(218));
F7219: entity F port map(lamdaA => P(7)(219),lamdaB => P(7)(223),lamdaOut => P(6)(219));
G7220: entity G port map(lamdaA => P(7)(216),lamdaB => P(7)(220),s => s(7)(108),lamdaOut => P(6)(220));
G7221: entity G port map(lamdaA => P(7)(217),lamdaB => P(7)(221),s => s(7)(109),lamdaOut => P(6)(221));
G7222: entity G port map(lamdaA => P(7)(218),lamdaB => P(7)(222),s => s(7)(110),lamdaOut => P(6)(222));
G7223: entity G port map(lamdaA => P(7)(219),lamdaB => P(7)(223),s => s(7)(111),lamdaOut => P(6)(223));
F7224: entity F port map(lamdaA => P(7)(224),lamdaB => P(7)(228),lamdaOut => P(6)(224));
F7225: entity F port map(lamdaA => P(7)(225),lamdaB => P(7)(229),lamdaOut => P(6)(225));
F7226: entity F port map(lamdaA => P(7)(226),lamdaB => P(7)(230),lamdaOut => P(6)(226));
F7227: entity F port map(lamdaA => P(7)(227),lamdaB => P(7)(231),lamdaOut => P(6)(227));
G7228: entity G port map(lamdaA => P(7)(224),lamdaB => P(7)(228),s => s(7)(112),lamdaOut => P(6)(228));
G7229: entity G port map(lamdaA => P(7)(225),lamdaB => P(7)(229),s => s(7)(113),lamdaOut => P(6)(229));
G7230: entity G port map(lamdaA => P(7)(226),lamdaB => P(7)(230),s => s(7)(114),lamdaOut => P(6)(230));
G7231: entity G port map(lamdaA => P(7)(227),lamdaB => P(7)(231),s => s(7)(115),lamdaOut => P(6)(231));
F7232: entity F port map(lamdaA => P(7)(232),lamdaB => P(7)(236),lamdaOut => P(6)(232));
F7233: entity F port map(lamdaA => P(7)(233),lamdaB => P(7)(237),lamdaOut => P(6)(233));
F7234: entity F port map(lamdaA => P(7)(234),lamdaB => P(7)(238),lamdaOut => P(6)(234));
F7235: entity F port map(lamdaA => P(7)(235),lamdaB => P(7)(239),lamdaOut => P(6)(235));
G7236: entity G port map(lamdaA => P(7)(232),lamdaB => P(7)(236),s => s(7)(116),lamdaOut => P(6)(236));
G7237: entity G port map(lamdaA => P(7)(233),lamdaB => P(7)(237),s => s(7)(117),lamdaOut => P(6)(237));
G7238: entity G port map(lamdaA => P(7)(234),lamdaB => P(7)(238),s => s(7)(118),lamdaOut => P(6)(238));
G7239: entity G port map(lamdaA => P(7)(235),lamdaB => P(7)(239),s => s(7)(119),lamdaOut => P(6)(239));
F7240: entity F port map(lamdaA => P(7)(240),lamdaB => P(7)(244),lamdaOut => P(6)(240));
F7241: entity F port map(lamdaA => P(7)(241),lamdaB => P(7)(245),lamdaOut => P(6)(241));
F7242: entity F port map(lamdaA => P(7)(242),lamdaB => P(7)(246),lamdaOut => P(6)(242));
F7243: entity F port map(lamdaA => P(7)(243),lamdaB => P(7)(247),lamdaOut => P(6)(243));
G7244: entity G port map(lamdaA => P(7)(240),lamdaB => P(7)(244),s => s(7)(120),lamdaOut => P(6)(244));
G7245: entity G port map(lamdaA => P(7)(241),lamdaB => P(7)(245),s => s(7)(121),lamdaOut => P(6)(245));
G7246: entity G port map(lamdaA => P(7)(242),lamdaB => P(7)(246),s => s(7)(122),lamdaOut => P(6)(246));
G7247: entity G port map(lamdaA => P(7)(243),lamdaB => P(7)(247),s => s(7)(123),lamdaOut => P(6)(247));
F7248: entity F port map(lamdaA => P(7)(248),lamdaB => P(7)(252),lamdaOut => P(6)(248));
F7249: entity F port map(lamdaA => P(7)(249),lamdaB => P(7)(253),lamdaOut => P(6)(249));
F7250: entity F port map(lamdaA => P(7)(250),lamdaB => P(7)(254),lamdaOut => P(6)(250));
F7251: entity F port map(lamdaA => P(7)(251),lamdaB => P(7)(255),lamdaOut => P(6)(251));
G7252: entity G port map(lamdaA => P(7)(248),lamdaB => P(7)(252),s => s(7)(124),lamdaOut => P(6)(252));
G7253: entity G port map(lamdaA => P(7)(249),lamdaB => P(7)(253),s => s(7)(125),lamdaOut => P(6)(253));
G7254: entity G port map(lamdaA => P(7)(250),lamdaB => P(7)(254),s => s(7)(126),lamdaOut => P(6)(254));
G7255: entity G port map(lamdaA => P(7)(251),lamdaB => P(7)(255),s => s(7)(127),lamdaOut => P(6)(255));
F7256: entity F port map(lamdaA => P(7)(256),lamdaB => P(7)(260),lamdaOut => P(6)(256));
F7257: entity F port map(lamdaA => P(7)(257),lamdaB => P(7)(261),lamdaOut => P(6)(257));
F7258: entity F port map(lamdaA => P(7)(258),lamdaB => P(7)(262),lamdaOut => P(6)(258));
F7259: entity F port map(lamdaA => P(7)(259),lamdaB => P(7)(263),lamdaOut => P(6)(259));
G7260: entity G port map(lamdaA => P(7)(256),lamdaB => P(7)(260),s => s(7)(128),lamdaOut => P(6)(260));
G7261: entity G port map(lamdaA => P(7)(257),lamdaB => P(7)(261),s => s(7)(129),lamdaOut => P(6)(261));
G7262: entity G port map(lamdaA => P(7)(258),lamdaB => P(7)(262),s => s(7)(130),lamdaOut => P(6)(262));
G7263: entity G port map(lamdaA => P(7)(259),lamdaB => P(7)(263),s => s(7)(131),lamdaOut => P(6)(263));
F7264: entity F port map(lamdaA => P(7)(264),lamdaB => P(7)(268),lamdaOut => P(6)(264));
F7265: entity F port map(lamdaA => P(7)(265),lamdaB => P(7)(269),lamdaOut => P(6)(265));
F7266: entity F port map(lamdaA => P(7)(266),lamdaB => P(7)(270),lamdaOut => P(6)(266));
F7267: entity F port map(lamdaA => P(7)(267),lamdaB => P(7)(271),lamdaOut => P(6)(267));
G7268: entity G port map(lamdaA => P(7)(264),lamdaB => P(7)(268),s => s(7)(132),lamdaOut => P(6)(268));
G7269: entity G port map(lamdaA => P(7)(265),lamdaB => P(7)(269),s => s(7)(133),lamdaOut => P(6)(269));
G7270: entity G port map(lamdaA => P(7)(266),lamdaB => P(7)(270),s => s(7)(134),lamdaOut => P(6)(270));
G7271: entity G port map(lamdaA => P(7)(267),lamdaB => P(7)(271),s => s(7)(135),lamdaOut => P(6)(271));
F7272: entity F port map(lamdaA => P(7)(272),lamdaB => P(7)(276),lamdaOut => P(6)(272));
F7273: entity F port map(lamdaA => P(7)(273),lamdaB => P(7)(277),lamdaOut => P(6)(273));
F7274: entity F port map(lamdaA => P(7)(274),lamdaB => P(7)(278),lamdaOut => P(6)(274));
F7275: entity F port map(lamdaA => P(7)(275),lamdaB => P(7)(279),lamdaOut => P(6)(275));
G7276: entity G port map(lamdaA => P(7)(272),lamdaB => P(7)(276),s => s(7)(136),lamdaOut => P(6)(276));
G7277: entity G port map(lamdaA => P(7)(273),lamdaB => P(7)(277),s => s(7)(137),lamdaOut => P(6)(277));
G7278: entity G port map(lamdaA => P(7)(274),lamdaB => P(7)(278),s => s(7)(138),lamdaOut => P(6)(278));
G7279: entity G port map(lamdaA => P(7)(275),lamdaB => P(7)(279),s => s(7)(139),lamdaOut => P(6)(279));
F7280: entity F port map(lamdaA => P(7)(280),lamdaB => P(7)(284),lamdaOut => P(6)(280));
F7281: entity F port map(lamdaA => P(7)(281),lamdaB => P(7)(285),lamdaOut => P(6)(281));
F7282: entity F port map(lamdaA => P(7)(282),lamdaB => P(7)(286),lamdaOut => P(6)(282));
F7283: entity F port map(lamdaA => P(7)(283),lamdaB => P(7)(287),lamdaOut => P(6)(283));
G7284: entity G port map(lamdaA => P(7)(280),lamdaB => P(7)(284),s => s(7)(140),lamdaOut => P(6)(284));
G7285: entity G port map(lamdaA => P(7)(281),lamdaB => P(7)(285),s => s(7)(141),lamdaOut => P(6)(285));
G7286: entity G port map(lamdaA => P(7)(282),lamdaB => P(7)(286),s => s(7)(142),lamdaOut => P(6)(286));
G7287: entity G port map(lamdaA => P(7)(283),lamdaB => P(7)(287),s => s(7)(143),lamdaOut => P(6)(287));
F7288: entity F port map(lamdaA => P(7)(288),lamdaB => P(7)(292),lamdaOut => P(6)(288));
F7289: entity F port map(lamdaA => P(7)(289),lamdaB => P(7)(293),lamdaOut => P(6)(289));
F7290: entity F port map(lamdaA => P(7)(290),lamdaB => P(7)(294),lamdaOut => P(6)(290));
F7291: entity F port map(lamdaA => P(7)(291),lamdaB => P(7)(295),lamdaOut => P(6)(291));
G7292: entity G port map(lamdaA => P(7)(288),lamdaB => P(7)(292),s => s(7)(144),lamdaOut => P(6)(292));
G7293: entity G port map(lamdaA => P(7)(289),lamdaB => P(7)(293),s => s(7)(145),lamdaOut => P(6)(293));
G7294: entity G port map(lamdaA => P(7)(290),lamdaB => P(7)(294),s => s(7)(146),lamdaOut => P(6)(294));
G7295: entity G port map(lamdaA => P(7)(291),lamdaB => P(7)(295),s => s(7)(147),lamdaOut => P(6)(295));
F7296: entity F port map(lamdaA => P(7)(296),lamdaB => P(7)(300),lamdaOut => P(6)(296));
F7297: entity F port map(lamdaA => P(7)(297),lamdaB => P(7)(301),lamdaOut => P(6)(297));
F7298: entity F port map(lamdaA => P(7)(298),lamdaB => P(7)(302),lamdaOut => P(6)(298));
F7299: entity F port map(lamdaA => P(7)(299),lamdaB => P(7)(303),lamdaOut => P(6)(299));
G7300: entity G port map(lamdaA => P(7)(296),lamdaB => P(7)(300),s => s(7)(148),lamdaOut => P(6)(300));
G7301: entity G port map(lamdaA => P(7)(297),lamdaB => P(7)(301),s => s(7)(149),lamdaOut => P(6)(301));
G7302: entity G port map(lamdaA => P(7)(298),lamdaB => P(7)(302),s => s(7)(150),lamdaOut => P(6)(302));
G7303: entity G port map(lamdaA => P(7)(299),lamdaB => P(7)(303),s => s(7)(151),lamdaOut => P(6)(303));
F7304: entity F port map(lamdaA => P(7)(304),lamdaB => P(7)(308),lamdaOut => P(6)(304));
F7305: entity F port map(lamdaA => P(7)(305),lamdaB => P(7)(309),lamdaOut => P(6)(305));
F7306: entity F port map(lamdaA => P(7)(306),lamdaB => P(7)(310),lamdaOut => P(6)(306));
F7307: entity F port map(lamdaA => P(7)(307),lamdaB => P(7)(311),lamdaOut => P(6)(307));
G7308: entity G port map(lamdaA => P(7)(304),lamdaB => P(7)(308),s => s(7)(152),lamdaOut => P(6)(308));
G7309: entity G port map(lamdaA => P(7)(305),lamdaB => P(7)(309),s => s(7)(153),lamdaOut => P(6)(309));
G7310: entity G port map(lamdaA => P(7)(306),lamdaB => P(7)(310),s => s(7)(154),lamdaOut => P(6)(310));
G7311: entity G port map(lamdaA => P(7)(307),lamdaB => P(7)(311),s => s(7)(155),lamdaOut => P(6)(311));
F7312: entity F port map(lamdaA => P(7)(312),lamdaB => P(7)(316),lamdaOut => P(6)(312));
F7313: entity F port map(lamdaA => P(7)(313),lamdaB => P(7)(317),lamdaOut => P(6)(313));
F7314: entity F port map(lamdaA => P(7)(314),lamdaB => P(7)(318),lamdaOut => P(6)(314));
F7315: entity F port map(lamdaA => P(7)(315),lamdaB => P(7)(319),lamdaOut => P(6)(315));
G7316: entity G port map(lamdaA => P(7)(312),lamdaB => P(7)(316),s => s(7)(156),lamdaOut => P(6)(316));
G7317: entity G port map(lamdaA => P(7)(313),lamdaB => P(7)(317),s => s(7)(157),lamdaOut => P(6)(317));
G7318: entity G port map(lamdaA => P(7)(314),lamdaB => P(7)(318),s => s(7)(158),lamdaOut => P(6)(318));
G7319: entity G port map(lamdaA => P(7)(315),lamdaB => P(7)(319),s => s(7)(159),lamdaOut => P(6)(319));
F7320: entity F port map(lamdaA => P(7)(320),lamdaB => P(7)(324),lamdaOut => P(6)(320));
F7321: entity F port map(lamdaA => P(7)(321),lamdaB => P(7)(325),lamdaOut => P(6)(321));
F7322: entity F port map(lamdaA => P(7)(322),lamdaB => P(7)(326),lamdaOut => P(6)(322));
F7323: entity F port map(lamdaA => P(7)(323),lamdaB => P(7)(327),lamdaOut => P(6)(323));
G7324: entity G port map(lamdaA => P(7)(320),lamdaB => P(7)(324),s => s(7)(160),lamdaOut => P(6)(324));
G7325: entity G port map(lamdaA => P(7)(321),lamdaB => P(7)(325),s => s(7)(161),lamdaOut => P(6)(325));
G7326: entity G port map(lamdaA => P(7)(322),lamdaB => P(7)(326),s => s(7)(162),lamdaOut => P(6)(326));
G7327: entity G port map(lamdaA => P(7)(323),lamdaB => P(7)(327),s => s(7)(163),lamdaOut => P(6)(327));
F7328: entity F port map(lamdaA => P(7)(328),lamdaB => P(7)(332),lamdaOut => P(6)(328));
F7329: entity F port map(lamdaA => P(7)(329),lamdaB => P(7)(333),lamdaOut => P(6)(329));
F7330: entity F port map(lamdaA => P(7)(330),lamdaB => P(7)(334),lamdaOut => P(6)(330));
F7331: entity F port map(lamdaA => P(7)(331),lamdaB => P(7)(335),lamdaOut => P(6)(331));
G7332: entity G port map(lamdaA => P(7)(328),lamdaB => P(7)(332),s => s(7)(164),lamdaOut => P(6)(332));
G7333: entity G port map(lamdaA => P(7)(329),lamdaB => P(7)(333),s => s(7)(165),lamdaOut => P(6)(333));
G7334: entity G port map(lamdaA => P(7)(330),lamdaB => P(7)(334),s => s(7)(166),lamdaOut => P(6)(334));
G7335: entity G port map(lamdaA => P(7)(331),lamdaB => P(7)(335),s => s(7)(167),lamdaOut => P(6)(335));
F7336: entity F port map(lamdaA => P(7)(336),lamdaB => P(7)(340),lamdaOut => P(6)(336));
F7337: entity F port map(lamdaA => P(7)(337),lamdaB => P(7)(341),lamdaOut => P(6)(337));
F7338: entity F port map(lamdaA => P(7)(338),lamdaB => P(7)(342),lamdaOut => P(6)(338));
F7339: entity F port map(lamdaA => P(7)(339),lamdaB => P(7)(343),lamdaOut => P(6)(339));
G7340: entity G port map(lamdaA => P(7)(336),lamdaB => P(7)(340),s => s(7)(168),lamdaOut => P(6)(340));
G7341: entity G port map(lamdaA => P(7)(337),lamdaB => P(7)(341),s => s(7)(169),lamdaOut => P(6)(341));
G7342: entity G port map(lamdaA => P(7)(338),lamdaB => P(7)(342),s => s(7)(170),lamdaOut => P(6)(342));
G7343: entity G port map(lamdaA => P(7)(339),lamdaB => P(7)(343),s => s(7)(171),lamdaOut => P(6)(343));
F7344: entity F port map(lamdaA => P(7)(344),lamdaB => P(7)(348),lamdaOut => P(6)(344));
F7345: entity F port map(lamdaA => P(7)(345),lamdaB => P(7)(349),lamdaOut => P(6)(345));
F7346: entity F port map(lamdaA => P(7)(346),lamdaB => P(7)(350),lamdaOut => P(6)(346));
F7347: entity F port map(lamdaA => P(7)(347),lamdaB => P(7)(351),lamdaOut => P(6)(347));
G7348: entity G port map(lamdaA => P(7)(344),lamdaB => P(7)(348),s => s(7)(172),lamdaOut => P(6)(348));
G7349: entity G port map(lamdaA => P(7)(345),lamdaB => P(7)(349),s => s(7)(173),lamdaOut => P(6)(349));
G7350: entity G port map(lamdaA => P(7)(346),lamdaB => P(7)(350),s => s(7)(174),lamdaOut => P(6)(350));
G7351: entity G port map(lamdaA => P(7)(347),lamdaB => P(7)(351),s => s(7)(175),lamdaOut => P(6)(351));
F7352: entity F port map(lamdaA => P(7)(352),lamdaB => P(7)(356),lamdaOut => P(6)(352));
F7353: entity F port map(lamdaA => P(7)(353),lamdaB => P(7)(357),lamdaOut => P(6)(353));
F7354: entity F port map(lamdaA => P(7)(354),lamdaB => P(7)(358),lamdaOut => P(6)(354));
F7355: entity F port map(lamdaA => P(7)(355),lamdaB => P(7)(359),lamdaOut => P(6)(355));
G7356: entity G port map(lamdaA => P(7)(352),lamdaB => P(7)(356),s => s(7)(176),lamdaOut => P(6)(356));
G7357: entity G port map(lamdaA => P(7)(353),lamdaB => P(7)(357),s => s(7)(177),lamdaOut => P(6)(357));
G7358: entity G port map(lamdaA => P(7)(354),lamdaB => P(7)(358),s => s(7)(178),lamdaOut => P(6)(358));
G7359: entity G port map(lamdaA => P(7)(355),lamdaB => P(7)(359),s => s(7)(179),lamdaOut => P(6)(359));
F7360: entity F port map(lamdaA => P(7)(360),lamdaB => P(7)(364),lamdaOut => P(6)(360));
F7361: entity F port map(lamdaA => P(7)(361),lamdaB => P(7)(365),lamdaOut => P(6)(361));
F7362: entity F port map(lamdaA => P(7)(362),lamdaB => P(7)(366),lamdaOut => P(6)(362));
F7363: entity F port map(lamdaA => P(7)(363),lamdaB => P(7)(367),lamdaOut => P(6)(363));
G7364: entity G port map(lamdaA => P(7)(360),lamdaB => P(7)(364),s => s(7)(180),lamdaOut => P(6)(364));
G7365: entity G port map(lamdaA => P(7)(361),lamdaB => P(7)(365),s => s(7)(181),lamdaOut => P(6)(365));
G7366: entity G port map(lamdaA => P(7)(362),lamdaB => P(7)(366),s => s(7)(182),lamdaOut => P(6)(366));
G7367: entity G port map(lamdaA => P(7)(363),lamdaB => P(7)(367),s => s(7)(183),lamdaOut => P(6)(367));
F7368: entity F port map(lamdaA => P(7)(368),lamdaB => P(7)(372),lamdaOut => P(6)(368));
F7369: entity F port map(lamdaA => P(7)(369),lamdaB => P(7)(373),lamdaOut => P(6)(369));
F7370: entity F port map(lamdaA => P(7)(370),lamdaB => P(7)(374),lamdaOut => P(6)(370));
F7371: entity F port map(lamdaA => P(7)(371),lamdaB => P(7)(375),lamdaOut => P(6)(371));
G7372: entity G port map(lamdaA => P(7)(368),lamdaB => P(7)(372),s => s(7)(184),lamdaOut => P(6)(372));
G7373: entity G port map(lamdaA => P(7)(369),lamdaB => P(7)(373),s => s(7)(185),lamdaOut => P(6)(373));
G7374: entity G port map(lamdaA => P(7)(370),lamdaB => P(7)(374),s => s(7)(186),lamdaOut => P(6)(374));
G7375: entity G port map(lamdaA => P(7)(371),lamdaB => P(7)(375),s => s(7)(187),lamdaOut => P(6)(375));
F7376: entity F port map(lamdaA => P(7)(376),lamdaB => P(7)(380),lamdaOut => P(6)(376));
F7377: entity F port map(lamdaA => P(7)(377),lamdaB => P(7)(381),lamdaOut => P(6)(377));
F7378: entity F port map(lamdaA => P(7)(378),lamdaB => P(7)(382),lamdaOut => P(6)(378));
F7379: entity F port map(lamdaA => P(7)(379),lamdaB => P(7)(383),lamdaOut => P(6)(379));
G7380: entity G port map(lamdaA => P(7)(376),lamdaB => P(7)(380),s => s(7)(188),lamdaOut => P(6)(380));
G7381: entity G port map(lamdaA => P(7)(377),lamdaB => P(7)(381),s => s(7)(189),lamdaOut => P(6)(381));
G7382: entity G port map(lamdaA => P(7)(378),lamdaB => P(7)(382),s => s(7)(190),lamdaOut => P(6)(382));
G7383: entity G port map(lamdaA => P(7)(379),lamdaB => P(7)(383),s => s(7)(191),lamdaOut => P(6)(383));
F7384: entity F port map(lamdaA => P(7)(384),lamdaB => P(7)(388),lamdaOut => P(6)(384));
F7385: entity F port map(lamdaA => P(7)(385),lamdaB => P(7)(389),lamdaOut => P(6)(385));
F7386: entity F port map(lamdaA => P(7)(386),lamdaB => P(7)(390),lamdaOut => P(6)(386));
F7387: entity F port map(lamdaA => P(7)(387),lamdaB => P(7)(391),lamdaOut => P(6)(387));
G7388: entity G port map(lamdaA => P(7)(384),lamdaB => P(7)(388),s => s(7)(192),lamdaOut => P(6)(388));
G7389: entity G port map(lamdaA => P(7)(385),lamdaB => P(7)(389),s => s(7)(193),lamdaOut => P(6)(389));
G7390: entity G port map(lamdaA => P(7)(386),lamdaB => P(7)(390),s => s(7)(194),lamdaOut => P(6)(390));
G7391: entity G port map(lamdaA => P(7)(387),lamdaB => P(7)(391),s => s(7)(195),lamdaOut => P(6)(391));
F7392: entity F port map(lamdaA => P(7)(392),lamdaB => P(7)(396),lamdaOut => P(6)(392));
F7393: entity F port map(lamdaA => P(7)(393),lamdaB => P(7)(397),lamdaOut => P(6)(393));
F7394: entity F port map(lamdaA => P(7)(394),lamdaB => P(7)(398),lamdaOut => P(6)(394));
F7395: entity F port map(lamdaA => P(7)(395),lamdaB => P(7)(399),lamdaOut => P(6)(395));
G7396: entity G port map(lamdaA => P(7)(392),lamdaB => P(7)(396),s => s(7)(196),lamdaOut => P(6)(396));
G7397: entity G port map(lamdaA => P(7)(393),lamdaB => P(7)(397),s => s(7)(197),lamdaOut => P(6)(397));
G7398: entity G port map(lamdaA => P(7)(394),lamdaB => P(7)(398),s => s(7)(198),lamdaOut => P(6)(398));
G7399: entity G port map(lamdaA => P(7)(395),lamdaB => P(7)(399),s => s(7)(199),lamdaOut => P(6)(399));
F7400: entity F port map(lamdaA => P(7)(400),lamdaB => P(7)(404),lamdaOut => P(6)(400));
F7401: entity F port map(lamdaA => P(7)(401),lamdaB => P(7)(405),lamdaOut => P(6)(401));
F7402: entity F port map(lamdaA => P(7)(402),lamdaB => P(7)(406),lamdaOut => P(6)(402));
F7403: entity F port map(lamdaA => P(7)(403),lamdaB => P(7)(407),lamdaOut => P(6)(403));
G7404: entity G port map(lamdaA => P(7)(400),lamdaB => P(7)(404),s => s(7)(200),lamdaOut => P(6)(404));
G7405: entity G port map(lamdaA => P(7)(401),lamdaB => P(7)(405),s => s(7)(201),lamdaOut => P(6)(405));
G7406: entity G port map(lamdaA => P(7)(402),lamdaB => P(7)(406),s => s(7)(202),lamdaOut => P(6)(406));
G7407: entity G port map(lamdaA => P(7)(403),lamdaB => P(7)(407),s => s(7)(203),lamdaOut => P(6)(407));
F7408: entity F port map(lamdaA => P(7)(408),lamdaB => P(7)(412),lamdaOut => P(6)(408));
F7409: entity F port map(lamdaA => P(7)(409),lamdaB => P(7)(413),lamdaOut => P(6)(409));
F7410: entity F port map(lamdaA => P(7)(410),lamdaB => P(7)(414),lamdaOut => P(6)(410));
F7411: entity F port map(lamdaA => P(7)(411),lamdaB => P(7)(415),lamdaOut => P(6)(411));
G7412: entity G port map(lamdaA => P(7)(408),lamdaB => P(7)(412),s => s(7)(204),lamdaOut => P(6)(412));
G7413: entity G port map(lamdaA => P(7)(409),lamdaB => P(7)(413),s => s(7)(205),lamdaOut => P(6)(413));
G7414: entity G port map(lamdaA => P(7)(410),lamdaB => P(7)(414),s => s(7)(206),lamdaOut => P(6)(414));
G7415: entity G port map(lamdaA => P(7)(411),lamdaB => P(7)(415),s => s(7)(207),lamdaOut => P(6)(415));
F7416: entity F port map(lamdaA => P(7)(416),lamdaB => P(7)(420),lamdaOut => P(6)(416));
F7417: entity F port map(lamdaA => P(7)(417),lamdaB => P(7)(421),lamdaOut => P(6)(417));
F7418: entity F port map(lamdaA => P(7)(418),lamdaB => P(7)(422),lamdaOut => P(6)(418));
F7419: entity F port map(lamdaA => P(7)(419),lamdaB => P(7)(423),lamdaOut => P(6)(419));
G7420: entity G port map(lamdaA => P(7)(416),lamdaB => P(7)(420),s => s(7)(208),lamdaOut => P(6)(420));
G7421: entity G port map(lamdaA => P(7)(417),lamdaB => P(7)(421),s => s(7)(209),lamdaOut => P(6)(421));
G7422: entity G port map(lamdaA => P(7)(418),lamdaB => P(7)(422),s => s(7)(210),lamdaOut => P(6)(422));
G7423: entity G port map(lamdaA => P(7)(419),lamdaB => P(7)(423),s => s(7)(211),lamdaOut => P(6)(423));
F7424: entity F port map(lamdaA => P(7)(424),lamdaB => P(7)(428),lamdaOut => P(6)(424));
F7425: entity F port map(lamdaA => P(7)(425),lamdaB => P(7)(429),lamdaOut => P(6)(425));
F7426: entity F port map(lamdaA => P(7)(426),lamdaB => P(7)(430),lamdaOut => P(6)(426));
F7427: entity F port map(lamdaA => P(7)(427),lamdaB => P(7)(431),lamdaOut => P(6)(427));
G7428: entity G port map(lamdaA => P(7)(424),lamdaB => P(7)(428),s => s(7)(212),lamdaOut => P(6)(428));
G7429: entity G port map(lamdaA => P(7)(425),lamdaB => P(7)(429),s => s(7)(213),lamdaOut => P(6)(429));
G7430: entity G port map(lamdaA => P(7)(426),lamdaB => P(7)(430),s => s(7)(214),lamdaOut => P(6)(430));
G7431: entity G port map(lamdaA => P(7)(427),lamdaB => P(7)(431),s => s(7)(215),lamdaOut => P(6)(431));
F7432: entity F port map(lamdaA => P(7)(432),lamdaB => P(7)(436),lamdaOut => P(6)(432));
F7433: entity F port map(lamdaA => P(7)(433),lamdaB => P(7)(437),lamdaOut => P(6)(433));
F7434: entity F port map(lamdaA => P(7)(434),lamdaB => P(7)(438),lamdaOut => P(6)(434));
F7435: entity F port map(lamdaA => P(7)(435),lamdaB => P(7)(439),lamdaOut => P(6)(435));
G7436: entity G port map(lamdaA => P(7)(432),lamdaB => P(7)(436),s => s(7)(216),lamdaOut => P(6)(436));
G7437: entity G port map(lamdaA => P(7)(433),lamdaB => P(7)(437),s => s(7)(217),lamdaOut => P(6)(437));
G7438: entity G port map(lamdaA => P(7)(434),lamdaB => P(7)(438),s => s(7)(218),lamdaOut => P(6)(438));
G7439: entity G port map(lamdaA => P(7)(435),lamdaB => P(7)(439),s => s(7)(219),lamdaOut => P(6)(439));
F7440: entity F port map(lamdaA => P(7)(440),lamdaB => P(7)(444),lamdaOut => P(6)(440));
F7441: entity F port map(lamdaA => P(7)(441),lamdaB => P(7)(445),lamdaOut => P(6)(441));
F7442: entity F port map(lamdaA => P(7)(442),lamdaB => P(7)(446),lamdaOut => P(6)(442));
F7443: entity F port map(lamdaA => P(7)(443),lamdaB => P(7)(447),lamdaOut => P(6)(443));
G7444: entity G port map(lamdaA => P(7)(440),lamdaB => P(7)(444),s => s(7)(220),lamdaOut => P(6)(444));
G7445: entity G port map(lamdaA => P(7)(441),lamdaB => P(7)(445),s => s(7)(221),lamdaOut => P(6)(445));
G7446: entity G port map(lamdaA => P(7)(442),lamdaB => P(7)(446),s => s(7)(222),lamdaOut => P(6)(446));
G7447: entity G port map(lamdaA => P(7)(443),lamdaB => P(7)(447),s => s(7)(223),lamdaOut => P(6)(447));
F7448: entity F port map(lamdaA => P(7)(448),lamdaB => P(7)(452),lamdaOut => P(6)(448));
F7449: entity F port map(lamdaA => P(7)(449),lamdaB => P(7)(453),lamdaOut => P(6)(449));
F7450: entity F port map(lamdaA => P(7)(450),lamdaB => P(7)(454),lamdaOut => P(6)(450));
F7451: entity F port map(lamdaA => P(7)(451),lamdaB => P(7)(455),lamdaOut => P(6)(451));
G7452: entity G port map(lamdaA => P(7)(448),lamdaB => P(7)(452),s => s(7)(224),lamdaOut => P(6)(452));
G7453: entity G port map(lamdaA => P(7)(449),lamdaB => P(7)(453),s => s(7)(225),lamdaOut => P(6)(453));
G7454: entity G port map(lamdaA => P(7)(450),lamdaB => P(7)(454),s => s(7)(226),lamdaOut => P(6)(454));
G7455: entity G port map(lamdaA => P(7)(451),lamdaB => P(7)(455),s => s(7)(227),lamdaOut => P(6)(455));
F7456: entity F port map(lamdaA => P(7)(456),lamdaB => P(7)(460),lamdaOut => P(6)(456));
F7457: entity F port map(lamdaA => P(7)(457),lamdaB => P(7)(461),lamdaOut => P(6)(457));
F7458: entity F port map(lamdaA => P(7)(458),lamdaB => P(7)(462),lamdaOut => P(6)(458));
F7459: entity F port map(lamdaA => P(7)(459),lamdaB => P(7)(463),lamdaOut => P(6)(459));
G7460: entity G port map(lamdaA => P(7)(456),lamdaB => P(7)(460),s => s(7)(228),lamdaOut => P(6)(460));
G7461: entity G port map(lamdaA => P(7)(457),lamdaB => P(7)(461),s => s(7)(229),lamdaOut => P(6)(461));
G7462: entity G port map(lamdaA => P(7)(458),lamdaB => P(7)(462),s => s(7)(230),lamdaOut => P(6)(462));
G7463: entity G port map(lamdaA => P(7)(459),lamdaB => P(7)(463),s => s(7)(231),lamdaOut => P(6)(463));
F7464: entity F port map(lamdaA => P(7)(464),lamdaB => P(7)(468),lamdaOut => P(6)(464));
F7465: entity F port map(lamdaA => P(7)(465),lamdaB => P(7)(469),lamdaOut => P(6)(465));
F7466: entity F port map(lamdaA => P(7)(466),lamdaB => P(7)(470),lamdaOut => P(6)(466));
F7467: entity F port map(lamdaA => P(7)(467),lamdaB => P(7)(471),lamdaOut => P(6)(467));
G7468: entity G port map(lamdaA => P(7)(464),lamdaB => P(7)(468),s => s(7)(232),lamdaOut => P(6)(468));
G7469: entity G port map(lamdaA => P(7)(465),lamdaB => P(7)(469),s => s(7)(233),lamdaOut => P(6)(469));
G7470: entity G port map(lamdaA => P(7)(466),lamdaB => P(7)(470),s => s(7)(234),lamdaOut => P(6)(470));
G7471: entity G port map(lamdaA => P(7)(467),lamdaB => P(7)(471),s => s(7)(235),lamdaOut => P(6)(471));
F7472: entity F port map(lamdaA => P(7)(472),lamdaB => P(7)(476),lamdaOut => P(6)(472));
F7473: entity F port map(lamdaA => P(7)(473),lamdaB => P(7)(477),lamdaOut => P(6)(473));
F7474: entity F port map(lamdaA => P(7)(474),lamdaB => P(7)(478),lamdaOut => P(6)(474));
F7475: entity F port map(lamdaA => P(7)(475),lamdaB => P(7)(479),lamdaOut => P(6)(475));
G7476: entity G port map(lamdaA => P(7)(472),lamdaB => P(7)(476),s => s(7)(236),lamdaOut => P(6)(476));
G7477: entity G port map(lamdaA => P(7)(473),lamdaB => P(7)(477),s => s(7)(237),lamdaOut => P(6)(477));
G7478: entity G port map(lamdaA => P(7)(474),lamdaB => P(7)(478),s => s(7)(238),lamdaOut => P(6)(478));
G7479: entity G port map(lamdaA => P(7)(475),lamdaB => P(7)(479),s => s(7)(239),lamdaOut => P(6)(479));
F7480: entity F port map(lamdaA => P(7)(480),lamdaB => P(7)(484),lamdaOut => P(6)(480));
F7481: entity F port map(lamdaA => P(7)(481),lamdaB => P(7)(485),lamdaOut => P(6)(481));
F7482: entity F port map(lamdaA => P(7)(482),lamdaB => P(7)(486),lamdaOut => P(6)(482));
F7483: entity F port map(lamdaA => P(7)(483),lamdaB => P(7)(487),lamdaOut => P(6)(483));
G7484: entity G port map(lamdaA => P(7)(480),lamdaB => P(7)(484),s => s(7)(240),lamdaOut => P(6)(484));
G7485: entity G port map(lamdaA => P(7)(481),lamdaB => P(7)(485),s => s(7)(241),lamdaOut => P(6)(485));
G7486: entity G port map(lamdaA => P(7)(482),lamdaB => P(7)(486),s => s(7)(242),lamdaOut => P(6)(486));
G7487: entity G port map(lamdaA => P(7)(483),lamdaB => P(7)(487),s => s(7)(243),lamdaOut => P(6)(487));
F7488: entity F port map(lamdaA => P(7)(488),lamdaB => P(7)(492),lamdaOut => P(6)(488));
F7489: entity F port map(lamdaA => P(7)(489),lamdaB => P(7)(493),lamdaOut => P(6)(489));
F7490: entity F port map(lamdaA => P(7)(490),lamdaB => P(7)(494),lamdaOut => P(6)(490));
F7491: entity F port map(lamdaA => P(7)(491),lamdaB => P(7)(495),lamdaOut => P(6)(491));
G7492: entity G port map(lamdaA => P(7)(488),lamdaB => P(7)(492),s => s(7)(244),lamdaOut => P(6)(492));
G7493: entity G port map(lamdaA => P(7)(489),lamdaB => P(7)(493),s => s(7)(245),lamdaOut => P(6)(493));
G7494: entity G port map(lamdaA => P(7)(490),lamdaB => P(7)(494),s => s(7)(246),lamdaOut => P(6)(494));
G7495: entity G port map(lamdaA => P(7)(491),lamdaB => P(7)(495),s => s(7)(247),lamdaOut => P(6)(495));
F7496: entity F port map(lamdaA => P(7)(496),lamdaB => P(7)(500),lamdaOut => P(6)(496));
F7497: entity F port map(lamdaA => P(7)(497),lamdaB => P(7)(501),lamdaOut => P(6)(497));
F7498: entity F port map(lamdaA => P(7)(498),lamdaB => P(7)(502),lamdaOut => P(6)(498));
F7499: entity F port map(lamdaA => P(7)(499),lamdaB => P(7)(503),lamdaOut => P(6)(499));
G7500: entity G port map(lamdaA => P(7)(496),lamdaB => P(7)(500),s => s(7)(248),lamdaOut => P(6)(500));
G7501: entity G port map(lamdaA => P(7)(497),lamdaB => P(7)(501),s => s(7)(249),lamdaOut => P(6)(501));
G7502: entity G port map(lamdaA => P(7)(498),lamdaB => P(7)(502),s => s(7)(250),lamdaOut => P(6)(502));
G7503: entity G port map(lamdaA => P(7)(499),lamdaB => P(7)(503),s => s(7)(251),lamdaOut => P(6)(503));
F7504: entity F port map(lamdaA => P(7)(504),lamdaB => P(7)(508),lamdaOut => P(6)(504));
F7505: entity F port map(lamdaA => P(7)(505),lamdaB => P(7)(509),lamdaOut => P(6)(505));
F7506: entity F port map(lamdaA => P(7)(506),lamdaB => P(7)(510),lamdaOut => P(6)(506));
F7507: entity F port map(lamdaA => P(7)(507),lamdaB => P(7)(511),lamdaOut => P(6)(507));
G7508: entity G port map(lamdaA => P(7)(504),lamdaB => P(7)(508),s => s(7)(252),lamdaOut => P(6)(508));
G7509: entity G port map(lamdaA => P(7)(505),lamdaB => P(7)(509),s => s(7)(253),lamdaOut => P(6)(509));
G7510: entity G port map(lamdaA => P(7)(506),lamdaB => P(7)(510),s => s(7)(254),lamdaOut => P(6)(510));
G7511: entity G port map(lamdaA => P(7)(507),lamdaB => P(7)(511),s => s(7)(255),lamdaOut => P(6)(511));
-- STAGE 6
F60: entity F port map(lamdaA => P(6)(0),lamdaB => P(6)(8),lamdaOut => P(5)(0));
F61: entity F port map(lamdaA => P(6)(1),lamdaB => P(6)(9),lamdaOut => P(5)(1));
F62: entity F port map(lamdaA => P(6)(2),lamdaB => P(6)(10),lamdaOut => P(5)(2));
F63: entity F port map(lamdaA => P(6)(3),lamdaB => P(6)(11),lamdaOut => P(5)(3));
F64: entity F port map(lamdaA => P(6)(4),lamdaB => P(6)(12),lamdaOut => P(5)(4));
F65: entity F port map(lamdaA => P(6)(5),lamdaB => P(6)(13),lamdaOut => P(5)(5));
F66: entity F port map(lamdaA => P(6)(6),lamdaB => P(6)(14),lamdaOut => P(5)(6));
F67: entity F port map(lamdaA => P(6)(7),lamdaB => P(6)(15),lamdaOut => P(5)(7));
G68: entity G port map(lamdaA => P(6)(0),lamdaB => P(6)(8),s => s(6)(0),lamdaOut => P(5)(8));
G69: entity G port map(lamdaA => P(6)(1),lamdaB => P(6)(9),s => s(6)(1),lamdaOut => P(5)(9));
G610: entity G port map(lamdaA => P(6)(2),lamdaB => P(6)(10),s => s(6)(2),lamdaOut => P(5)(10));
G611: entity G port map(lamdaA => P(6)(3),lamdaB => P(6)(11),s => s(6)(3),lamdaOut => P(5)(11));
G612: entity G port map(lamdaA => P(6)(4),lamdaB => P(6)(12),s => s(6)(4),lamdaOut => P(5)(12));
G613: entity G port map(lamdaA => P(6)(5),lamdaB => P(6)(13),s => s(6)(5),lamdaOut => P(5)(13));
G614: entity G port map(lamdaA => P(6)(6),lamdaB => P(6)(14),s => s(6)(6),lamdaOut => P(5)(14));
G615: entity G port map(lamdaA => P(6)(7),lamdaB => P(6)(15),s => s(6)(7),lamdaOut => P(5)(15));
F616: entity F port map(lamdaA => P(6)(16),lamdaB => P(6)(24),lamdaOut => P(5)(16));
F617: entity F port map(lamdaA => P(6)(17),lamdaB => P(6)(25),lamdaOut => P(5)(17));
F618: entity F port map(lamdaA => P(6)(18),lamdaB => P(6)(26),lamdaOut => P(5)(18));
F619: entity F port map(lamdaA => P(6)(19),lamdaB => P(6)(27),lamdaOut => P(5)(19));
F620: entity F port map(lamdaA => P(6)(20),lamdaB => P(6)(28),lamdaOut => P(5)(20));
F621: entity F port map(lamdaA => P(6)(21),lamdaB => P(6)(29),lamdaOut => P(5)(21));
F622: entity F port map(lamdaA => P(6)(22),lamdaB => P(6)(30),lamdaOut => P(5)(22));
F623: entity F port map(lamdaA => P(6)(23),lamdaB => P(6)(31),lamdaOut => P(5)(23));
G624: entity G port map(lamdaA => P(6)(16),lamdaB => P(6)(24),s => s(6)(8),lamdaOut => P(5)(24));
G625: entity G port map(lamdaA => P(6)(17),lamdaB => P(6)(25),s => s(6)(9),lamdaOut => P(5)(25));
G626: entity G port map(lamdaA => P(6)(18),lamdaB => P(6)(26),s => s(6)(10),lamdaOut => P(5)(26));
G627: entity G port map(lamdaA => P(6)(19),lamdaB => P(6)(27),s => s(6)(11),lamdaOut => P(5)(27));
G628: entity G port map(lamdaA => P(6)(20),lamdaB => P(6)(28),s => s(6)(12),lamdaOut => P(5)(28));
G629: entity G port map(lamdaA => P(6)(21),lamdaB => P(6)(29),s => s(6)(13),lamdaOut => P(5)(29));
G630: entity G port map(lamdaA => P(6)(22),lamdaB => P(6)(30),s => s(6)(14),lamdaOut => P(5)(30));
G631: entity G port map(lamdaA => P(6)(23),lamdaB => P(6)(31),s => s(6)(15),lamdaOut => P(5)(31));
F632: entity F port map(lamdaA => P(6)(32),lamdaB => P(6)(40),lamdaOut => P(5)(32));
F633: entity F port map(lamdaA => P(6)(33),lamdaB => P(6)(41),lamdaOut => P(5)(33));
F634: entity F port map(lamdaA => P(6)(34),lamdaB => P(6)(42),lamdaOut => P(5)(34));
F635: entity F port map(lamdaA => P(6)(35),lamdaB => P(6)(43),lamdaOut => P(5)(35));
F636: entity F port map(lamdaA => P(6)(36),lamdaB => P(6)(44),lamdaOut => P(5)(36));
F637: entity F port map(lamdaA => P(6)(37),lamdaB => P(6)(45),lamdaOut => P(5)(37));
F638: entity F port map(lamdaA => P(6)(38),lamdaB => P(6)(46),lamdaOut => P(5)(38));
F639: entity F port map(lamdaA => P(6)(39),lamdaB => P(6)(47),lamdaOut => P(5)(39));
G640: entity G port map(lamdaA => P(6)(32),lamdaB => P(6)(40),s => s(6)(16),lamdaOut => P(5)(40));
G641: entity G port map(lamdaA => P(6)(33),lamdaB => P(6)(41),s => s(6)(17),lamdaOut => P(5)(41));
G642: entity G port map(lamdaA => P(6)(34),lamdaB => P(6)(42),s => s(6)(18),lamdaOut => P(5)(42));
G643: entity G port map(lamdaA => P(6)(35),lamdaB => P(6)(43),s => s(6)(19),lamdaOut => P(5)(43));
G644: entity G port map(lamdaA => P(6)(36),lamdaB => P(6)(44),s => s(6)(20),lamdaOut => P(5)(44));
G645: entity G port map(lamdaA => P(6)(37),lamdaB => P(6)(45),s => s(6)(21),lamdaOut => P(5)(45));
G646: entity G port map(lamdaA => P(6)(38),lamdaB => P(6)(46),s => s(6)(22),lamdaOut => P(5)(46));
G647: entity G port map(lamdaA => P(6)(39),lamdaB => P(6)(47),s => s(6)(23),lamdaOut => P(5)(47));
F648: entity F port map(lamdaA => P(6)(48),lamdaB => P(6)(56),lamdaOut => P(5)(48));
F649: entity F port map(lamdaA => P(6)(49),lamdaB => P(6)(57),lamdaOut => P(5)(49));
F650: entity F port map(lamdaA => P(6)(50),lamdaB => P(6)(58),lamdaOut => P(5)(50));
F651: entity F port map(lamdaA => P(6)(51),lamdaB => P(6)(59),lamdaOut => P(5)(51));
F652: entity F port map(lamdaA => P(6)(52),lamdaB => P(6)(60),lamdaOut => P(5)(52));
F653: entity F port map(lamdaA => P(6)(53),lamdaB => P(6)(61),lamdaOut => P(5)(53));
F654: entity F port map(lamdaA => P(6)(54),lamdaB => P(6)(62),lamdaOut => P(5)(54));
F655: entity F port map(lamdaA => P(6)(55),lamdaB => P(6)(63),lamdaOut => P(5)(55));
G656: entity G port map(lamdaA => P(6)(48),lamdaB => P(6)(56),s => s(6)(24),lamdaOut => P(5)(56));
G657: entity G port map(lamdaA => P(6)(49),lamdaB => P(6)(57),s => s(6)(25),lamdaOut => P(5)(57));
G658: entity G port map(lamdaA => P(6)(50),lamdaB => P(6)(58),s => s(6)(26),lamdaOut => P(5)(58));
G659: entity G port map(lamdaA => P(6)(51),lamdaB => P(6)(59),s => s(6)(27),lamdaOut => P(5)(59));
G660: entity G port map(lamdaA => P(6)(52),lamdaB => P(6)(60),s => s(6)(28),lamdaOut => P(5)(60));
G661: entity G port map(lamdaA => P(6)(53),lamdaB => P(6)(61),s => s(6)(29),lamdaOut => P(5)(61));
G662: entity G port map(lamdaA => P(6)(54),lamdaB => P(6)(62),s => s(6)(30),lamdaOut => P(5)(62));
G663: entity G port map(lamdaA => P(6)(55),lamdaB => P(6)(63),s => s(6)(31),lamdaOut => P(5)(63));
F664: entity F port map(lamdaA => P(6)(64),lamdaB => P(6)(72),lamdaOut => P(5)(64));
F665: entity F port map(lamdaA => P(6)(65),lamdaB => P(6)(73),lamdaOut => P(5)(65));
F666: entity F port map(lamdaA => P(6)(66),lamdaB => P(6)(74),lamdaOut => P(5)(66));
F667: entity F port map(lamdaA => P(6)(67),lamdaB => P(6)(75),lamdaOut => P(5)(67));
F668: entity F port map(lamdaA => P(6)(68),lamdaB => P(6)(76),lamdaOut => P(5)(68));
F669: entity F port map(lamdaA => P(6)(69),lamdaB => P(6)(77),lamdaOut => P(5)(69));
F670: entity F port map(lamdaA => P(6)(70),lamdaB => P(6)(78),lamdaOut => P(5)(70));
F671: entity F port map(lamdaA => P(6)(71),lamdaB => P(6)(79),lamdaOut => P(5)(71));
G672: entity G port map(lamdaA => P(6)(64),lamdaB => P(6)(72),s => s(6)(32),lamdaOut => P(5)(72));
G673: entity G port map(lamdaA => P(6)(65),lamdaB => P(6)(73),s => s(6)(33),lamdaOut => P(5)(73));
G674: entity G port map(lamdaA => P(6)(66),lamdaB => P(6)(74),s => s(6)(34),lamdaOut => P(5)(74));
G675: entity G port map(lamdaA => P(6)(67),lamdaB => P(6)(75),s => s(6)(35),lamdaOut => P(5)(75));
G676: entity G port map(lamdaA => P(6)(68),lamdaB => P(6)(76),s => s(6)(36),lamdaOut => P(5)(76));
G677: entity G port map(lamdaA => P(6)(69),lamdaB => P(6)(77),s => s(6)(37),lamdaOut => P(5)(77));
G678: entity G port map(lamdaA => P(6)(70),lamdaB => P(6)(78),s => s(6)(38),lamdaOut => P(5)(78));
G679: entity G port map(lamdaA => P(6)(71),lamdaB => P(6)(79),s => s(6)(39),lamdaOut => P(5)(79));
F680: entity F port map(lamdaA => P(6)(80),lamdaB => P(6)(88),lamdaOut => P(5)(80));
F681: entity F port map(lamdaA => P(6)(81),lamdaB => P(6)(89),lamdaOut => P(5)(81));
F682: entity F port map(lamdaA => P(6)(82),lamdaB => P(6)(90),lamdaOut => P(5)(82));
F683: entity F port map(lamdaA => P(6)(83),lamdaB => P(6)(91),lamdaOut => P(5)(83));
F684: entity F port map(lamdaA => P(6)(84),lamdaB => P(6)(92),lamdaOut => P(5)(84));
F685: entity F port map(lamdaA => P(6)(85),lamdaB => P(6)(93),lamdaOut => P(5)(85));
F686: entity F port map(lamdaA => P(6)(86),lamdaB => P(6)(94),lamdaOut => P(5)(86));
F687: entity F port map(lamdaA => P(6)(87),lamdaB => P(6)(95),lamdaOut => P(5)(87));
G688: entity G port map(lamdaA => P(6)(80),lamdaB => P(6)(88),s => s(6)(40),lamdaOut => P(5)(88));
G689: entity G port map(lamdaA => P(6)(81),lamdaB => P(6)(89),s => s(6)(41),lamdaOut => P(5)(89));
G690: entity G port map(lamdaA => P(6)(82),lamdaB => P(6)(90),s => s(6)(42),lamdaOut => P(5)(90));
G691: entity G port map(lamdaA => P(6)(83),lamdaB => P(6)(91),s => s(6)(43),lamdaOut => P(5)(91));
G692: entity G port map(lamdaA => P(6)(84),lamdaB => P(6)(92),s => s(6)(44),lamdaOut => P(5)(92));
G693: entity G port map(lamdaA => P(6)(85),lamdaB => P(6)(93),s => s(6)(45),lamdaOut => P(5)(93));
G694: entity G port map(lamdaA => P(6)(86),lamdaB => P(6)(94),s => s(6)(46),lamdaOut => P(5)(94));
G695: entity G port map(lamdaA => P(6)(87),lamdaB => P(6)(95),s => s(6)(47),lamdaOut => P(5)(95));
F696: entity F port map(lamdaA => P(6)(96),lamdaB => P(6)(104),lamdaOut => P(5)(96));
F697: entity F port map(lamdaA => P(6)(97),lamdaB => P(6)(105),lamdaOut => P(5)(97));
F698: entity F port map(lamdaA => P(6)(98),lamdaB => P(6)(106),lamdaOut => P(5)(98));
F699: entity F port map(lamdaA => P(6)(99),lamdaB => P(6)(107),lamdaOut => P(5)(99));
F6100: entity F port map(lamdaA => P(6)(100),lamdaB => P(6)(108),lamdaOut => P(5)(100));
F6101: entity F port map(lamdaA => P(6)(101),lamdaB => P(6)(109),lamdaOut => P(5)(101));
F6102: entity F port map(lamdaA => P(6)(102),lamdaB => P(6)(110),lamdaOut => P(5)(102));
F6103: entity F port map(lamdaA => P(6)(103),lamdaB => P(6)(111),lamdaOut => P(5)(103));
G6104: entity G port map(lamdaA => P(6)(96),lamdaB => P(6)(104),s => s(6)(48),lamdaOut => P(5)(104));
G6105: entity G port map(lamdaA => P(6)(97),lamdaB => P(6)(105),s => s(6)(49),lamdaOut => P(5)(105));
G6106: entity G port map(lamdaA => P(6)(98),lamdaB => P(6)(106),s => s(6)(50),lamdaOut => P(5)(106));
G6107: entity G port map(lamdaA => P(6)(99),lamdaB => P(6)(107),s => s(6)(51),lamdaOut => P(5)(107));
G6108: entity G port map(lamdaA => P(6)(100),lamdaB => P(6)(108),s => s(6)(52),lamdaOut => P(5)(108));
G6109: entity G port map(lamdaA => P(6)(101),lamdaB => P(6)(109),s => s(6)(53),lamdaOut => P(5)(109));
G6110: entity G port map(lamdaA => P(6)(102),lamdaB => P(6)(110),s => s(6)(54),lamdaOut => P(5)(110));
G6111: entity G port map(lamdaA => P(6)(103),lamdaB => P(6)(111),s => s(6)(55),lamdaOut => P(5)(111));
F6112: entity F port map(lamdaA => P(6)(112),lamdaB => P(6)(120),lamdaOut => P(5)(112));
F6113: entity F port map(lamdaA => P(6)(113),lamdaB => P(6)(121),lamdaOut => P(5)(113));
F6114: entity F port map(lamdaA => P(6)(114),lamdaB => P(6)(122),lamdaOut => P(5)(114));
F6115: entity F port map(lamdaA => P(6)(115),lamdaB => P(6)(123),lamdaOut => P(5)(115));
F6116: entity F port map(lamdaA => P(6)(116),lamdaB => P(6)(124),lamdaOut => P(5)(116));
F6117: entity F port map(lamdaA => P(6)(117),lamdaB => P(6)(125),lamdaOut => P(5)(117));
F6118: entity F port map(lamdaA => P(6)(118),lamdaB => P(6)(126),lamdaOut => P(5)(118));
F6119: entity F port map(lamdaA => P(6)(119),lamdaB => P(6)(127),lamdaOut => P(5)(119));
G6120: entity G port map(lamdaA => P(6)(112),lamdaB => P(6)(120),s => s(6)(56),lamdaOut => P(5)(120));
G6121: entity G port map(lamdaA => P(6)(113),lamdaB => P(6)(121),s => s(6)(57),lamdaOut => P(5)(121));
G6122: entity G port map(lamdaA => P(6)(114),lamdaB => P(6)(122),s => s(6)(58),lamdaOut => P(5)(122));
G6123: entity G port map(lamdaA => P(6)(115),lamdaB => P(6)(123),s => s(6)(59),lamdaOut => P(5)(123));
G6124: entity G port map(lamdaA => P(6)(116),lamdaB => P(6)(124),s => s(6)(60),lamdaOut => P(5)(124));
G6125: entity G port map(lamdaA => P(6)(117),lamdaB => P(6)(125),s => s(6)(61),lamdaOut => P(5)(125));
G6126: entity G port map(lamdaA => P(6)(118),lamdaB => P(6)(126),s => s(6)(62),lamdaOut => P(5)(126));
G6127: entity G port map(lamdaA => P(6)(119),lamdaB => P(6)(127),s => s(6)(63),lamdaOut => P(5)(127));
F6128: entity F port map(lamdaA => P(6)(128),lamdaB => P(6)(136),lamdaOut => P(5)(128));
F6129: entity F port map(lamdaA => P(6)(129),lamdaB => P(6)(137),lamdaOut => P(5)(129));
F6130: entity F port map(lamdaA => P(6)(130),lamdaB => P(6)(138),lamdaOut => P(5)(130));
F6131: entity F port map(lamdaA => P(6)(131),lamdaB => P(6)(139),lamdaOut => P(5)(131));
F6132: entity F port map(lamdaA => P(6)(132),lamdaB => P(6)(140),lamdaOut => P(5)(132));
F6133: entity F port map(lamdaA => P(6)(133),lamdaB => P(6)(141),lamdaOut => P(5)(133));
F6134: entity F port map(lamdaA => P(6)(134),lamdaB => P(6)(142),lamdaOut => P(5)(134));
F6135: entity F port map(lamdaA => P(6)(135),lamdaB => P(6)(143),lamdaOut => P(5)(135));
G6136: entity G port map(lamdaA => P(6)(128),lamdaB => P(6)(136),s => s(6)(64),lamdaOut => P(5)(136));
G6137: entity G port map(lamdaA => P(6)(129),lamdaB => P(6)(137),s => s(6)(65),lamdaOut => P(5)(137));
G6138: entity G port map(lamdaA => P(6)(130),lamdaB => P(6)(138),s => s(6)(66),lamdaOut => P(5)(138));
G6139: entity G port map(lamdaA => P(6)(131),lamdaB => P(6)(139),s => s(6)(67),lamdaOut => P(5)(139));
G6140: entity G port map(lamdaA => P(6)(132),lamdaB => P(6)(140),s => s(6)(68),lamdaOut => P(5)(140));
G6141: entity G port map(lamdaA => P(6)(133),lamdaB => P(6)(141),s => s(6)(69),lamdaOut => P(5)(141));
G6142: entity G port map(lamdaA => P(6)(134),lamdaB => P(6)(142),s => s(6)(70),lamdaOut => P(5)(142));
G6143: entity G port map(lamdaA => P(6)(135),lamdaB => P(6)(143),s => s(6)(71),lamdaOut => P(5)(143));
F6144: entity F port map(lamdaA => P(6)(144),lamdaB => P(6)(152),lamdaOut => P(5)(144));
F6145: entity F port map(lamdaA => P(6)(145),lamdaB => P(6)(153),lamdaOut => P(5)(145));
F6146: entity F port map(lamdaA => P(6)(146),lamdaB => P(6)(154),lamdaOut => P(5)(146));
F6147: entity F port map(lamdaA => P(6)(147),lamdaB => P(6)(155),lamdaOut => P(5)(147));
F6148: entity F port map(lamdaA => P(6)(148),lamdaB => P(6)(156),lamdaOut => P(5)(148));
F6149: entity F port map(lamdaA => P(6)(149),lamdaB => P(6)(157),lamdaOut => P(5)(149));
F6150: entity F port map(lamdaA => P(6)(150),lamdaB => P(6)(158),lamdaOut => P(5)(150));
F6151: entity F port map(lamdaA => P(6)(151),lamdaB => P(6)(159),lamdaOut => P(5)(151));
G6152: entity G port map(lamdaA => P(6)(144),lamdaB => P(6)(152),s => s(6)(72),lamdaOut => P(5)(152));
G6153: entity G port map(lamdaA => P(6)(145),lamdaB => P(6)(153),s => s(6)(73),lamdaOut => P(5)(153));
G6154: entity G port map(lamdaA => P(6)(146),lamdaB => P(6)(154),s => s(6)(74),lamdaOut => P(5)(154));
G6155: entity G port map(lamdaA => P(6)(147),lamdaB => P(6)(155),s => s(6)(75),lamdaOut => P(5)(155));
G6156: entity G port map(lamdaA => P(6)(148),lamdaB => P(6)(156),s => s(6)(76),lamdaOut => P(5)(156));
G6157: entity G port map(lamdaA => P(6)(149),lamdaB => P(6)(157),s => s(6)(77),lamdaOut => P(5)(157));
G6158: entity G port map(lamdaA => P(6)(150),lamdaB => P(6)(158),s => s(6)(78),lamdaOut => P(5)(158));
G6159: entity G port map(lamdaA => P(6)(151),lamdaB => P(6)(159),s => s(6)(79),lamdaOut => P(5)(159));
F6160: entity F port map(lamdaA => P(6)(160),lamdaB => P(6)(168),lamdaOut => P(5)(160));
F6161: entity F port map(lamdaA => P(6)(161),lamdaB => P(6)(169),lamdaOut => P(5)(161));
F6162: entity F port map(lamdaA => P(6)(162),lamdaB => P(6)(170),lamdaOut => P(5)(162));
F6163: entity F port map(lamdaA => P(6)(163),lamdaB => P(6)(171),lamdaOut => P(5)(163));
F6164: entity F port map(lamdaA => P(6)(164),lamdaB => P(6)(172),lamdaOut => P(5)(164));
F6165: entity F port map(lamdaA => P(6)(165),lamdaB => P(6)(173),lamdaOut => P(5)(165));
F6166: entity F port map(lamdaA => P(6)(166),lamdaB => P(6)(174),lamdaOut => P(5)(166));
F6167: entity F port map(lamdaA => P(6)(167),lamdaB => P(6)(175),lamdaOut => P(5)(167));
G6168: entity G port map(lamdaA => P(6)(160),lamdaB => P(6)(168),s => s(6)(80),lamdaOut => P(5)(168));
G6169: entity G port map(lamdaA => P(6)(161),lamdaB => P(6)(169),s => s(6)(81),lamdaOut => P(5)(169));
G6170: entity G port map(lamdaA => P(6)(162),lamdaB => P(6)(170),s => s(6)(82),lamdaOut => P(5)(170));
G6171: entity G port map(lamdaA => P(6)(163),lamdaB => P(6)(171),s => s(6)(83),lamdaOut => P(5)(171));
G6172: entity G port map(lamdaA => P(6)(164),lamdaB => P(6)(172),s => s(6)(84),lamdaOut => P(5)(172));
G6173: entity G port map(lamdaA => P(6)(165),lamdaB => P(6)(173),s => s(6)(85),lamdaOut => P(5)(173));
G6174: entity G port map(lamdaA => P(6)(166),lamdaB => P(6)(174),s => s(6)(86),lamdaOut => P(5)(174));
G6175: entity G port map(lamdaA => P(6)(167),lamdaB => P(6)(175),s => s(6)(87),lamdaOut => P(5)(175));
F6176: entity F port map(lamdaA => P(6)(176),lamdaB => P(6)(184),lamdaOut => P(5)(176));
F6177: entity F port map(lamdaA => P(6)(177),lamdaB => P(6)(185),lamdaOut => P(5)(177));
F6178: entity F port map(lamdaA => P(6)(178),lamdaB => P(6)(186),lamdaOut => P(5)(178));
F6179: entity F port map(lamdaA => P(6)(179),lamdaB => P(6)(187),lamdaOut => P(5)(179));
F6180: entity F port map(lamdaA => P(6)(180),lamdaB => P(6)(188),lamdaOut => P(5)(180));
F6181: entity F port map(lamdaA => P(6)(181),lamdaB => P(6)(189),lamdaOut => P(5)(181));
F6182: entity F port map(lamdaA => P(6)(182),lamdaB => P(6)(190),lamdaOut => P(5)(182));
F6183: entity F port map(lamdaA => P(6)(183),lamdaB => P(6)(191),lamdaOut => P(5)(183));
G6184: entity G port map(lamdaA => P(6)(176),lamdaB => P(6)(184),s => s(6)(88),lamdaOut => P(5)(184));
G6185: entity G port map(lamdaA => P(6)(177),lamdaB => P(6)(185),s => s(6)(89),lamdaOut => P(5)(185));
G6186: entity G port map(lamdaA => P(6)(178),lamdaB => P(6)(186),s => s(6)(90),lamdaOut => P(5)(186));
G6187: entity G port map(lamdaA => P(6)(179),lamdaB => P(6)(187),s => s(6)(91),lamdaOut => P(5)(187));
G6188: entity G port map(lamdaA => P(6)(180),lamdaB => P(6)(188),s => s(6)(92),lamdaOut => P(5)(188));
G6189: entity G port map(lamdaA => P(6)(181),lamdaB => P(6)(189),s => s(6)(93),lamdaOut => P(5)(189));
G6190: entity G port map(lamdaA => P(6)(182),lamdaB => P(6)(190),s => s(6)(94),lamdaOut => P(5)(190));
G6191: entity G port map(lamdaA => P(6)(183),lamdaB => P(6)(191),s => s(6)(95),lamdaOut => P(5)(191));
F6192: entity F port map(lamdaA => P(6)(192),lamdaB => P(6)(200),lamdaOut => P(5)(192));
F6193: entity F port map(lamdaA => P(6)(193),lamdaB => P(6)(201),lamdaOut => P(5)(193));
F6194: entity F port map(lamdaA => P(6)(194),lamdaB => P(6)(202),lamdaOut => P(5)(194));
F6195: entity F port map(lamdaA => P(6)(195),lamdaB => P(6)(203),lamdaOut => P(5)(195));
F6196: entity F port map(lamdaA => P(6)(196),lamdaB => P(6)(204),lamdaOut => P(5)(196));
F6197: entity F port map(lamdaA => P(6)(197),lamdaB => P(6)(205),lamdaOut => P(5)(197));
F6198: entity F port map(lamdaA => P(6)(198),lamdaB => P(6)(206),lamdaOut => P(5)(198));
F6199: entity F port map(lamdaA => P(6)(199),lamdaB => P(6)(207),lamdaOut => P(5)(199));
G6200: entity G port map(lamdaA => P(6)(192),lamdaB => P(6)(200),s => s(6)(96),lamdaOut => P(5)(200));
G6201: entity G port map(lamdaA => P(6)(193),lamdaB => P(6)(201),s => s(6)(97),lamdaOut => P(5)(201));
G6202: entity G port map(lamdaA => P(6)(194),lamdaB => P(6)(202),s => s(6)(98),lamdaOut => P(5)(202));
G6203: entity G port map(lamdaA => P(6)(195),lamdaB => P(6)(203),s => s(6)(99),lamdaOut => P(5)(203));
G6204: entity G port map(lamdaA => P(6)(196),lamdaB => P(6)(204),s => s(6)(100),lamdaOut => P(5)(204));
G6205: entity G port map(lamdaA => P(6)(197),lamdaB => P(6)(205),s => s(6)(101),lamdaOut => P(5)(205));
G6206: entity G port map(lamdaA => P(6)(198),lamdaB => P(6)(206),s => s(6)(102),lamdaOut => P(5)(206));
G6207: entity G port map(lamdaA => P(6)(199),lamdaB => P(6)(207),s => s(6)(103),lamdaOut => P(5)(207));
F6208: entity F port map(lamdaA => P(6)(208),lamdaB => P(6)(216),lamdaOut => P(5)(208));
F6209: entity F port map(lamdaA => P(6)(209),lamdaB => P(6)(217),lamdaOut => P(5)(209));
F6210: entity F port map(lamdaA => P(6)(210),lamdaB => P(6)(218),lamdaOut => P(5)(210));
F6211: entity F port map(lamdaA => P(6)(211),lamdaB => P(6)(219),lamdaOut => P(5)(211));
F6212: entity F port map(lamdaA => P(6)(212),lamdaB => P(6)(220),lamdaOut => P(5)(212));
F6213: entity F port map(lamdaA => P(6)(213),lamdaB => P(6)(221),lamdaOut => P(5)(213));
F6214: entity F port map(lamdaA => P(6)(214),lamdaB => P(6)(222),lamdaOut => P(5)(214));
F6215: entity F port map(lamdaA => P(6)(215),lamdaB => P(6)(223),lamdaOut => P(5)(215));
G6216: entity G port map(lamdaA => P(6)(208),lamdaB => P(6)(216),s => s(6)(104),lamdaOut => P(5)(216));
G6217: entity G port map(lamdaA => P(6)(209),lamdaB => P(6)(217),s => s(6)(105),lamdaOut => P(5)(217));
G6218: entity G port map(lamdaA => P(6)(210),lamdaB => P(6)(218),s => s(6)(106),lamdaOut => P(5)(218));
G6219: entity G port map(lamdaA => P(6)(211),lamdaB => P(6)(219),s => s(6)(107),lamdaOut => P(5)(219));
G6220: entity G port map(lamdaA => P(6)(212),lamdaB => P(6)(220),s => s(6)(108),lamdaOut => P(5)(220));
G6221: entity G port map(lamdaA => P(6)(213),lamdaB => P(6)(221),s => s(6)(109),lamdaOut => P(5)(221));
G6222: entity G port map(lamdaA => P(6)(214),lamdaB => P(6)(222),s => s(6)(110),lamdaOut => P(5)(222));
G6223: entity G port map(lamdaA => P(6)(215),lamdaB => P(6)(223),s => s(6)(111),lamdaOut => P(5)(223));
F6224: entity F port map(lamdaA => P(6)(224),lamdaB => P(6)(232),lamdaOut => P(5)(224));
F6225: entity F port map(lamdaA => P(6)(225),lamdaB => P(6)(233),lamdaOut => P(5)(225));
F6226: entity F port map(lamdaA => P(6)(226),lamdaB => P(6)(234),lamdaOut => P(5)(226));
F6227: entity F port map(lamdaA => P(6)(227),lamdaB => P(6)(235),lamdaOut => P(5)(227));
F6228: entity F port map(lamdaA => P(6)(228),lamdaB => P(6)(236),lamdaOut => P(5)(228));
F6229: entity F port map(lamdaA => P(6)(229),lamdaB => P(6)(237),lamdaOut => P(5)(229));
F6230: entity F port map(lamdaA => P(6)(230),lamdaB => P(6)(238),lamdaOut => P(5)(230));
F6231: entity F port map(lamdaA => P(6)(231),lamdaB => P(6)(239),lamdaOut => P(5)(231));
G6232: entity G port map(lamdaA => P(6)(224),lamdaB => P(6)(232),s => s(6)(112),lamdaOut => P(5)(232));
G6233: entity G port map(lamdaA => P(6)(225),lamdaB => P(6)(233),s => s(6)(113),lamdaOut => P(5)(233));
G6234: entity G port map(lamdaA => P(6)(226),lamdaB => P(6)(234),s => s(6)(114),lamdaOut => P(5)(234));
G6235: entity G port map(lamdaA => P(6)(227),lamdaB => P(6)(235),s => s(6)(115),lamdaOut => P(5)(235));
G6236: entity G port map(lamdaA => P(6)(228),lamdaB => P(6)(236),s => s(6)(116),lamdaOut => P(5)(236));
G6237: entity G port map(lamdaA => P(6)(229),lamdaB => P(6)(237),s => s(6)(117),lamdaOut => P(5)(237));
G6238: entity G port map(lamdaA => P(6)(230),lamdaB => P(6)(238),s => s(6)(118),lamdaOut => P(5)(238));
G6239: entity G port map(lamdaA => P(6)(231),lamdaB => P(6)(239),s => s(6)(119),lamdaOut => P(5)(239));
F6240: entity F port map(lamdaA => P(6)(240),lamdaB => P(6)(248),lamdaOut => P(5)(240));
F6241: entity F port map(lamdaA => P(6)(241),lamdaB => P(6)(249),lamdaOut => P(5)(241));
F6242: entity F port map(lamdaA => P(6)(242),lamdaB => P(6)(250),lamdaOut => P(5)(242));
F6243: entity F port map(lamdaA => P(6)(243),lamdaB => P(6)(251),lamdaOut => P(5)(243));
F6244: entity F port map(lamdaA => P(6)(244),lamdaB => P(6)(252),lamdaOut => P(5)(244));
F6245: entity F port map(lamdaA => P(6)(245),lamdaB => P(6)(253),lamdaOut => P(5)(245));
F6246: entity F port map(lamdaA => P(6)(246),lamdaB => P(6)(254),lamdaOut => P(5)(246));
F6247: entity F port map(lamdaA => P(6)(247),lamdaB => P(6)(255),lamdaOut => P(5)(247));
G6248: entity G port map(lamdaA => P(6)(240),lamdaB => P(6)(248),s => s(6)(120),lamdaOut => P(5)(248));
G6249: entity G port map(lamdaA => P(6)(241),lamdaB => P(6)(249),s => s(6)(121),lamdaOut => P(5)(249));
G6250: entity G port map(lamdaA => P(6)(242),lamdaB => P(6)(250),s => s(6)(122),lamdaOut => P(5)(250));
G6251: entity G port map(lamdaA => P(6)(243),lamdaB => P(6)(251),s => s(6)(123),lamdaOut => P(5)(251));
G6252: entity G port map(lamdaA => P(6)(244),lamdaB => P(6)(252),s => s(6)(124),lamdaOut => P(5)(252));
G6253: entity G port map(lamdaA => P(6)(245),lamdaB => P(6)(253),s => s(6)(125),lamdaOut => P(5)(253));
G6254: entity G port map(lamdaA => P(6)(246),lamdaB => P(6)(254),s => s(6)(126),lamdaOut => P(5)(254));
G6255: entity G port map(lamdaA => P(6)(247),lamdaB => P(6)(255),s => s(6)(127),lamdaOut => P(5)(255));
F6256: entity F port map(lamdaA => P(6)(256),lamdaB => P(6)(264),lamdaOut => P(5)(256));
F6257: entity F port map(lamdaA => P(6)(257),lamdaB => P(6)(265),lamdaOut => P(5)(257));
F6258: entity F port map(lamdaA => P(6)(258),lamdaB => P(6)(266),lamdaOut => P(5)(258));
F6259: entity F port map(lamdaA => P(6)(259),lamdaB => P(6)(267),lamdaOut => P(5)(259));
F6260: entity F port map(lamdaA => P(6)(260),lamdaB => P(6)(268),lamdaOut => P(5)(260));
F6261: entity F port map(lamdaA => P(6)(261),lamdaB => P(6)(269),lamdaOut => P(5)(261));
F6262: entity F port map(lamdaA => P(6)(262),lamdaB => P(6)(270),lamdaOut => P(5)(262));
F6263: entity F port map(lamdaA => P(6)(263),lamdaB => P(6)(271),lamdaOut => P(5)(263));
G6264: entity G port map(lamdaA => P(6)(256),lamdaB => P(6)(264),s => s(6)(128),lamdaOut => P(5)(264));
G6265: entity G port map(lamdaA => P(6)(257),lamdaB => P(6)(265),s => s(6)(129),lamdaOut => P(5)(265));
G6266: entity G port map(lamdaA => P(6)(258),lamdaB => P(6)(266),s => s(6)(130),lamdaOut => P(5)(266));
G6267: entity G port map(lamdaA => P(6)(259),lamdaB => P(6)(267),s => s(6)(131),lamdaOut => P(5)(267));
G6268: entity G port map(lamdaA => P(6)(260),lamdaB => P(6)(268),s => s(6)(132),lamdaOut => P(5)(268));
G6269: entity G port map(lamdaA => P(6)(261),lamdaB => P(6)(269),s => s(6)(133),lamdaOut => P(5)(269));
G6270: entity G port map(lamdaA => P(6)(262),lamdaB => P(6)(270),s => s(6)(134),lamdaOut => P(5)(270));
G6271: entity G port map(lamdaA => P(6)(263),lamdaB => P(6)(271),s => s(6)(135),lamdaOut => P(5)(271));
F6272: entity F port map(lamdaA => P(6)(272),lamdaB => P(6)(280),lamdaOut => P(5)(272));
F6273: entity F port map(lamdaA => P(6)(273),lamdaB => P(6)(281),lamdaOut => P(5)(273));
F6274: entity F port map(lamdaA => P(6)(274),lamdaB => P(6)(282),lamdaOut => P(5)(274));
F6275: entity F port map(lamdaA => P(6)(275),lamdaB => P(6)(283),lamdaOut => P(5)(275));
F6276: entity F port map(lamdaA => P(6)(276),lamdaB => P(6)(284),lamdaOut => P(5)(276));
F6277: entity F port map(lamdaA => P(6)(277),lamdaB => P(6)(285),lamdaOut => P(5)(277));
F6278: entity F port map(lamdaA => P(6)(278),lamdaB => P(6)(286),lamdaOut => P(5)(278));
F6279: entity F port map(lamdaA => P(6)(279),lamdaB => P(6)(287),lamdaOut => P(5)(279));
G6280: entity G port map(lamdaA => P(6)(272),lamdaB => P(6)(280),s => s(6)(136),lamdaOut => P(5)(280));
G6281: entity G port map(lamdaA => P(6)(273),lamdaB => P(6)(281),s => s(6)(137),lamdaOut => P(5)(281));
G6282: entity G port map(lamdaA => P(6)(274),lamdaB => P(6)(282),s => s(6)(138),lamdaOut => P(5)(282));
G6283: entity G port map(lamdaA => P(6)(275),lamdaB => P(6)(283),s => s(6)(139),lamdaOut => P(5)(283));
G6284: entity G port map(lamdaA => P(6)(276),lamdaB => P(6)(284),s => s(6)(140),lamdaOut => P(5)(284));
G6285: entity G port map(lamdaA => P(6)(277),lamdaB => P(6)(285),s => s(6)(141),lamdaOut => P(5)(285));
G6286: entity G port map(lamdaA => P(6)(278),lamdaB => P(6)(286),s => s(6)(142),lamdaOut => P(5)(286));
G6287: entity G port map(lamdaA => P(6)(279),lamdaB => P(6)(287),s => s(6)(143),lamdaOut => P(5)(287));
F6288: entity F port map(lamdaA => P(6)(288),lamdaB => P(6)(296),lamdaOut => P(5)(288));
F6289: entity F port map(lamdaA => P(6)(289),lamdaB => P(6)(297),lamdaOut => P(5)(289));
F6290: entity F port map(lamdaA => P(6)(290),lamdaB => P(6)(298),lamdaOut => P(5)(290));
F6291: entity F port map(lamdaA => P(6)(291),lamdaB => P(6)(299),lamdaOut => P(5)(291));
F6292: entity F port map(lamdaA => P(6)(292),lamdaB => P(6)(300),lamdaOut => P(5)(292));
F6293: entity F port map(lamdaA => P(6)(293),lamdaB => P(6)(301),lamdaOut => P(5)(293));
F6294: entity F port map(lamdaA => P(6)(294),lamdaB => P(6)(302),lamdaOut => P(5)(294));
F6295: entity F port map(lamdaA => P(6)(295),lamdaB => P(6)(303),lamdaOut => P(5)(295));
G6296: entity G port map(lamdaA => P(6)(288),lamdaB => P(6)(296),s => s(6)(144),lamdaOut => P(5)(296));
G6297: entity G port map(lamdaA => P(6)(289),lamdaB => P(6)(297),s => s(6)(145),lamdaOut => P(5)(297));
G6298: entity G port map(lamdaA => P(6)(290),lamdaB => P(6)(298),s => s(6)(146),lamdaOut => P(5)(298));
G6299: entity G port map(lamdaA => P(6)(291),lamdaB => P(6)(299),s => s(6)(147),lamdaOut => P(5)(299));
G6300: entity G port map(lamdaA => P(6)(292),lamdaB => P(6)(300),s => s(6)(148),lamdaOut => P(5)(300));
G6301: entity G port map(lamdaA => P(6)(293),lamdaB => P(6)(301),s => s(6)(149),lamdaOut => P(5)(301));
G6302: entity G port map(lamdaA => P(6)(294),lamdaB => P(6)(302),s => s(6)(150),lamdaOut => P(5)(302));
G6303: entity G port map(lamdaA => P(6)(295),lamdaB => P(6)(303),s => s(6)(151),lamdaOut => P(5)(303));
F6304: entity F port map(lamdaA => P(6)(304),lamdaB => P(6)(312),lamdaOut => P(5)(304));
F6305: entity F port map(lamdaA => P(6)(305),lamdaB => P(6)(313),lamdaOut => P(5)(305));
F6306: entity F port map(lamdaA => P(6)(306),lamdaB => P(6)(314),lamdaOut => P(5)(306));
F6307: entity F port map(lamdaA => P(6)(307),lamdaB => P(6)(315),lamdaOut => P(5)(307));
F6308: entity F port map(lamdaA => P(6)(308),lamdaB => P(6)(316),lamdaOut => P(5)(308));
F6309: entity F port map(lamdaA => P(6)(309),lamdaB => P(6)(317),lamdaOut => P(5)(309));
F6310: entity F port map(lamdaA => P(6)(310),lamdaB => P(6)(318),lamdaOut => P(5)(310));
F6311: entity F port map(lamdaA => P(6)(311),lamdaB => P(6)(319),lamdaOut => P(5)(311));
G6312: entity G port map(lamdaA => P(6)(304),lamdaB => P(6)(312),s => s(6)(152),lamdaOut => P(5)(312));
G6313: entity G port map(lamdaA => P(6)(305),lamdaB => P(6)(313),s => s(6)(153),lamdaOut => P(5)(313));
G6314: entity G port map(lamdaA => P(6)(306),lamdaB => P(6)(314),s => s(6)(154),lamdaOut => P(5)(314));
G6315: entity G port map(lamdaA => P(6)(307),lamdaB => P(6)(315),s => s(6)(155),lamdaOut => P(5)(315));
G6316: entity G port map(lamdaA => P(6)(308),lamdaB => P(6)(316),s => s(6)(156),lamdaOut => P(5)(316));
G6317: entity G port map(lamdaA => P(6)(309),lamdaB => P(6)(317),s => s(6)(157),lamdaOut => P(5)(317));
G6318: entity G port map(lamdaA => P(6)(310),lamdaB => P(6)(318),s => s(6)(158),lamdaOut => P(5)(318));
G6319: entity G port map(lamdaA => P(6)(311),lamdaB => P(6)(319),s => s(6)(159),lamdaOut => P(5)(319));
F6320: entity F port map(lamdaA => P(6)(320),lamdaB => P(6)(328),lamdaOut => P(5)(320));
F6321: entity F port map(lamdaA => P(6)(321),lamdaB => P(6)(329),lamdaOut => P(5)(321));
F6322: entity F port map(lamdaA => P(6)(322),lamdaB => P(6)(330),lamdaOut => P(5)(322));
F6323: entity F port map(lamdaA => P(6)(323),lamdaB => P(6)(331),lamdaOut => P(5)(323));
F6324: entity F port map(lamdaA => P(6)(324),lamdaB => P(6)(332),lamdaOut => P(5)(324));
F6325: entity F port map(lamdaA => P(6)(325),lamdaB => P(6)(333),lamdaOut => P(5)(325));
F6326: entity F port map(lamdaA => P(6)(326),lamdaB => P(6)(334),lamdaOut => P(5)(326));
F6327: entity F port map(lamdaA => P(6)(327),lamdaB => P(6)(335),lamdaOut => P(5)(327));
G6328: entity G port map(lamdaA => P(6)(320),lamdaB => P(6)(328),s => s(6)(160),lamdaOut => P(5)(328));
G6329: entity G port map(lamdaA => P(6)(321),lamdaB => P(6)(329),s => s(6)(161),lamdaOut => P(5)(329));
G6330: entity G port map(lamdaA => P(6)(322),lamdaB => P(6)(330),s => s(6)(162),lamdaOut => P(5)(330));
G6331: entity G port map(lamdaA => P(6)(323),lamdaB => P(6)(331),s => s(6)(163),lamdaOut => P(5)(331));
G6332: entity G port map(lamdaA => P(6)(324),lamdaB => P(6)(332),s => s(6)(164),lamdaOut => P(5)(332));
G6333: entity G port map(lamdaA => P(6)(325),lamdaB => P(6)(333),s => s(6)(165),lamdaOut => P(5)(333));
G6334: entity G port map(lamdaA => P(6)(326),lamdaB => P(6)(334),s => s(6)(166),lamdaOut => P(5)(334));
G6335: entity G port map(lamdaA => P(6)(327),lamdaB => P(6)(335),s => s(6)(167),lamdaOut => P(5)(335));
F6336: entity F port map(lamdaA => P(6)(336),lamdaB => P(6)(344),lamdaOut => P(5)(336));
F6337: entity F port map(lamdaA => P(6)(337),lamdaB => P(6)(345),lamdaOut => P(5)(337));
F6338: entity F port map(lamdaA => P(6)(338),lamdaB => P(6)(346),lamdaOut => P(5)(338));
F6339: entity F port map(lamdaA => P(6)(339),lamdaB => P(6)(347),lamdaOut => P(5)(339));
F6340: entity F port map(lamdaA => P(6)(340),lamdaB => P(6)(348),lamdaOut => P(5)(340));
F6341: entity F port map(lamdaA => P(6)(341),lamdaB => P(6)(349),lamdaOut => P(5)(341));
F6342: entity F port map(lamdaA => P(6)(342),lamdaB => P(6)(350),lamdaOut => P(5)(342));
F6343: entity F port map(lamdaA => P(6)(343),lamdaB => P(6)(351),lamdaOut => P(5)(343));
G6344: entity G port map(lamdaA => P(6)(336),lamdaB => P(6)(344),s => s(6)(168),lamdaOut => P(5)(344));
G6345: entity G port map(lamdaA => P(6)(337),lamdaB => P(6)(345),s => s(6)(169),lamdaOut => P(5)(345));
G6346: entity G port map(lamdaA => P(6)(338),lamdaB => P(6)(346),s => s(6)(170),lamdaOut => P(5)(346));
G6347: entity G port map(lamdaA => P(6)(339),lamdaB => P(6)(347),s => s(6)(171),lamdaOut => P(5)(347));
G6348: entity G port map(lamdaA => P(6)(340),lamdaB => P(6)(348),s => s(6)(172),lamdaOut => P(5)(348));
G6349: entity G port map(lamdaA => P(6)(341),lamdaB => P(6)(349),s => s(6)(173),lamdaOut => P(5)(349));
G6350: entity G port map(lamdaA => P(6)(342),lamdaB => P(6)(350),s => s(6)(174),lamdaOut => P(5)(350));
G6351: entity G port map(lamdaA => P(6)(343),lamdaB => P(6)(351),s => s(6)(175),lamdaOut => P(5)(351));
F6352: entity F port map(lamdaA => P(6)(352),lamdaB => P(6)(360),lamdaOut => P(5)(352));
F6353: entity F port map(lamdaA => P(6)(353),lamdaB => P(6)(361),lamdaOut => P(5)(353));
F6354: entity F port map(lamdaA => P(6)(354),lamdaB => P(6)(362),lamdaOut => P(5)(354));
F6355: entity F port map(lamdaA => P(6)(355),lamdaB => P(6)(363),lamdaOut => P(5)(355));
F6356: entity F port map(lamdaA => P(6)(356),lamdaB => P(6)(364),lamdaOut => P(5)(356));
F6357: entity F port map(lamdaA => P(6)(357),lamdaB => P(6)(365),lamdaOut => P(5)(357));
F6358: entity F port map(lamdaA => P(6)(358),lamdaB => P(6)(366),lamdaOut => P(5)(358));
F6359: entity F port map(lamdaA => P(6)(359),lamdaB => P(6)(367),lamdaOut => P(5)(359));
G6360: entity G port map(lamdaA => P(6)(352),lamdaB => P(6)(360),s => s(6)(176),lamdaOut => P(5)(360));
G6361: entity G port map(lamdaA => P(6)(353),lamdaB => P(6)(361),s => s(6)(177),lamdaOut => P(5)(361));
G6362: entity G port map(lamdaA => P(6)(354),lamdaB => P(6)(362),s => s(6)(178),lamdaOut => P(5)(362));
G6363: entity G port map(lamdaA => P(6)(355),lamdaB => P(6)(363),s => s(6)(179),lamdaOut => P(5)(363));
G6364: entity G port map(lamdaA => P(6)(356),lamdaB => P(6)(364),s => s(6)(180),lamdaOut => P(5)(364));
G6365: entity G port map(lamdaA => P(6)(357),lamdaB => P(6)(365),s => s(6)(181),lamdaOut => P(5)(365));
G6366: entity G port map(lamdaA => P(6)(358),lamdaB => P(6)(366),s => s(6)(182),lamdaOut => P(5)(366));
G6367: entity G port map(lamdaA => P(6)(359),lamdaB => P(6)(367),s => s(6)(183),lamdaOut => P(5)(367));
F6368: entity F port map(lamdaA => P(6)(368),lamdaB => P(6)(376),lamdaOut => P(5)(368));
F6369: entity F port map(lamdaA => P(6)(369),lamdaB => P(6)(377),lamdaOut => P(5)(369));
F6370: entity F port map(lamdaA => P(6)(370),lamdaB => P(6)(378),lamdaOut => P(5)(370));
F6371: entity F port map(lamdaA => P(6)(371),lamdaB => P(6)(379),lamdaOut => P(5)(371));
F6372: entity F port map(lamdaA => P(6)(372),lamdaB => P(6)(380),lamdaOut => P(5)(372));
F6373: entity F port map(lamdaA => P(6)(373),lamdaB => P(6)(381),lamdaOut => P(5)(373));
F6374: entity F port map(lamdaA => P(6)(374),lamdaB => P(6)(382),lamdaOut => P(5)(374));
F6375: entity F port map(lamdaA => P(6)(375),lamdaB => P(6)(383),lamdaOut => P(5)(375));
G6376: entity G port map(lamdaA => P(6)(368),lamdaB => P(6)(376),s => s(6)(184),lamdaOut => P(5)(376));
G6377: entity G port map(lamdaA => P(6)(369),lamdaB => P(6)(377),s => s(6)(185),lamdaOut => P(5)(377));
G6378: entity G port map(lamdaA => P(6)(370),lamdaB => P(6)(378),s => s(6)(186),lamdaOut => P(5)(378));
G6379: entity G port map(lamdaA => P(6)(371),lamdaB => P(6)(379),s => s(6)(187),lamdaOut => P(5)(379));
G6380: entity G port map(lamdaA => P(6)(372),lamdaB => P(6)(380),s => s(6)(188),lamdaOut => P(5)(380));
G6381: entity G port map(lamdaA => P(6)(373),lamdaB => P(6)(381),s => s(6)(189),lamdaOut => P(5)(381));
G6382: entity G port map(lamdaA => P(6)(374),lamdaB => P(6)(382),s => s(6)(190),lamdaOut => P(5)(382));
G6383: entity G port map(lamdaA => P(6)(375),lamdaB => P(6)(383),s => s(6)(191),lamdaOut => P(5)(383));
F6384: entity F port map(lamdaA => P(6)(384),lamdaB => P(6)(392),lamdaOut => P(5)(384));
F6385: entity F port map(lamdaA => P(6)(385),lamdaB => P(6)(393),lamdaOut => P(5)(385));
F6386: entity F port map(lamdaA => P(6)(386),lamdaB => P(6)(394),lamdaOut => P(5)(386));
F6387: entity F port map(lamdaA => P(6)(387),lamdaB => P(6)(395),lamdaOut => P(5)(387));
F6388: entity F port map(lamdaA => P(6)(388),lamdaB => P(6)(396),lamdaOut => P(5)(388));
F6389: entity F port map(lamdaA => P(6)(389),lamdaB => P(6)(397),lamdaOut => P(5)(389));
F6390: entity F port map(lamdaA => P(6)(390),lamdaB => P(6)(398),lamdaOut => P(5)(390));
F6391: entity F port map(lamdaA => P(6)(391),lamdaB => P(6)(399),lamdaOut => P(5)(391));
G6392: entity G port map(lamdaA => P(6)(384),lamdaB => P(6)(392),s => s(6)(192),lamdaOut => P(5)(392));
G6393: entity G port map(lamdaA => P(6)(385),lamdaB => P(6)(393),s => s(6)(193),lamdaOut => P(5)(393));
G6394: entity G port map(lamdaA => P(6)(386),lamdaB => P(6)(394),s => s(6)(194),lamdaOut => P(5)(394));
G6395: entity G port map(lamdaA => P(6)(387),lamdaB => P(6)(395),s => s(6)(195),lamdaOut => P(5)(395));
G6396: entity G port map(lamdaA => P(6)(388),lamdaB => P(6)(396),s => s(6)(196),lamdaOut => P(5)(396));
G6397: entity G port map(lamdaA => P(6)(389),lamdaB => P(6)(397),s => s(6)(197),lamdaOut => P(5)(397));
G6398: entity G port map(lamdaA => P(6)(390),lamdaB => P(6)(398),s => s(6)(198),lamdaOut => P(5)(398));
G6399: entity G port map(lamdaA => P(6)(391),lamdaB => P(6)(399),s => s(6)(199),lamdaOut => P(5)(399));
F6400: entity F port map(lamdaA => P(6)(400),lamdaB => P(6)(408),lamdaOut => P(5)(400));
F6401: entity F port map(lamdaA => P(6)(401),lamdaB => P(6)(409),lamdaOut => P(5)(401));
F6402: entity F port map(lamdaA => P(6)(402),lamdaB => P(6)(410),lamdaOut => P(5)(402));
F6403: entity F port map(lamdaA => P(6)(403),lamdaB => P(6)(411),lamdaOut => P(5)(403));
F6404: entity F port map(lamdaA => P(6)(404),lamdaB => P(6)(412),lamdaOut => P(5)(404));
F6405: entity F port map(lamdaA => P(6)(405),lamdaB => P(6)(413),lamdaOut => P(5)(405));
F6406: entity F port map(lamdaA => P(6)(406),lamdaB => P(6)(414),lamdaOut => P(5)(406));
F6407: entity F port map(lamdaA => P(6)(407),lamdaB => P(6)(415),lamdaOut => P(5)(407));
G6408: entity G port map(lamdaA => P(6)(400),lamdaB => P(6)(408),s => s(6)(200),lamdaOut => P(5)(408));
G6409: entity G port map(lamdaA => P(6)(401),lamdaB => P(6)(409),s => s(6)(201),lamdaOut => P(5)(409));
G6410: entity G port map(lamdaA => P(6)(402),lamdaB => P(6)(410),s => s(6)(202),lamdaOut => P(5)(410));
G6411: entity G port map(lamdaA => P(6)(403),lamdaB => P(6)(411),s => s(6)(203),lamdaOut => P(5)(411));
G6412: entity G port map(lamdaA => P(6)(404),lamdaB => P(6)(412),s => s(6)(204),lamdaOut => P(5)(412));
G6413: entity G port map(lamdaA => P(6)(405),lamdaB => P(6)(413),s => s(6)(205),lamdaOut => P(5)(413));
G6414: entity G port map(lamdaA => P(6)(406),lamdaB => P(6)(414),s => s(6)(206),lamdaOut => P(5)(414));
G6415: entity G port map(lamdaA => P(6)(407),lamdaB => P(6)(415),s => s(6)(207),lamdaOut => P(5)(415));
F6416: entity F port map(lamdaA => P(6)(416),lamdaB => P(6)(424),lamdaOut => P(5)(416));
F6417: entity F port map(lamdaA => P(6)(417),lamdaB => P(6)(425),lamdaOut => P(5)(417));
F6418: entity F port map(lamdaA => P(6)(418),lamdaB => P(6)(426),lamdaOut => P(5)(418));
F6419: entity F port map(lamdaA => P(6)(419),lamdaB => P(6)(427),lamdaOut => P(5)(419));
F6420: entity F port map(lamdaA => P(6)(420),lamdaB => P(6)(428),lamdaOut => P(5)(420));
F6421: entity F port map(lamdaA => P(6)(421),lamdaB => P(6)(429),lamdaOut => P(5)(421));
F6422: entity F port map(lamdaA => P(6)(422),lamdaB => P(6)(430),lamdaOut => P(5)(422));
F6423: entity F port map(lamdaA => P(6)(423),lamdaB => P(6)(431),lamdaOut => P(5)(423));
G6424: entity G port map(lamdaA => P(6)(416),lamdaB => P(6)(424),s => s(6)(208),lamdaOut => P(5)(424));
G6425: entity G port map(lamdaA => P(6)(417),lamdaB => P(6)(425),s => s(6)(209),lamdaOut => P(5)(425));
G6426: entity G port map(lamdaA => P(6)(418),lamdaB => P(6)(426),s => s(6)(210),lamdaOut => P(5)(426));
G6427: entity G port map(lamdaA => P(6)(419),lamdaB => P(6)(427),s => s(6)(211),lamdaOut => P(5)(427));
G6428: entity G port map(lamdaA => P(6)(420),lamdaB => P(6)(428),s => s(6)(212),lamdaOut => P(5)(428));
G6429: entity G port map(lamdaA => P(6)(421),lamdaB => P(6)(429),s => s(6)(213),lamdaOut => P(5)(429));
G6430: entity G port map(lamdaA => P(6)(422),lamdaB => P(6)(430),s => s(6)(214),lamdaOut => P(5)(430));
G6431: entity G port map(lamdaA => P(6)(423),lamdaB => P(6)(431),s => s(6)(215),lamdaOut => P(5)(431));
F6432: entity F port map(lamdaA => P(6)(432),lamdaB => P(6)(440),lamdaOut => P(5)(432));
F6433: entity F port map(lamdaA => P(6)(433),lamdaB => P(6)(441),lamdaOut => P(5)(433));
F6434: entity F port map(lamdaA => P(6)(434),lamdaB => P(6)(442),lamdaOut => P(5)(434));
F6435: entity F port map(lamdaA => P(6)(435),lamdaB => P(6)(443),lamdaOut => P(5)(435));
F6436: entity F port map(lamdaA => P(6)(436),lamdaB => P(6)(444),lamdaOut => P(5)(436));
F6437: entity F port map(lamdaA => P(6)(437),lamdaB => P(6)(445),lamdaOut => P(5)(437));
F6438: entity F port map(lamdaA => P(6)(438),lamdaB => P(6)(446),lamdaOut => P(5)(438));
F6439: entity F port map(lamdaA => P(6)(439),lamdaB => P(6)(447),lamdaOut => P(5)(439));
G6440: entity G port map(lamdaA => P(6)(432),lamdaB => P(6)(440),s => s(6)(216),lamdaOut => P(5)(440));
G6441: entity G port map(lamdaA => P(6)(433),lamdaB => P(6)(441),s => s(6)(217),lamdaOut => P(5)(441));
G6442: entity G port map(lamdaA => P(6)(434),lamdaB => P(6)(442),s => s(6)(218),lamdaOut => P(5)(442));
G6443: entity G port map(lamdaA => P(6)(435),lamdaB => P(6)(443),s => s(6)(219),lamdaOut => P(5)(443));
G6444: entity G port map(lamdaA => P(6)(436),lamdaB => P(6)(444),s => s(6)(220),lamdaOut => P(5)(444));
G6445: entity G port map(lamdaA => P(6)(437),lamdaB => P(6)(445),s => s(6)(221),lamdaOut => P(5)(445));
G6446: entity G port map(lamdaA => P(6)(438),lamdaB => P(6)(446),s => s(6)(222),lamdaOut => P(5)(446));
G6447: entity G port map(lamdaA => P(6)(439),lamdaB => P(6)(447),s => s(6)(223),lamdaOut => P(5)(447));
F6448: entity F port map(lamdaA => P(6)(448),lamdaB => P(6)(456),lamdaOut => P(5)(448));
F6449: entity F port map(lamdaA => P(6)(449),lamdaB => P(6)(457),lamdaOut => P(5)(449));
F6450: entity F port map(lamdaA => P(6)(450),lamdaB => P(6)(458),lamdaOut => P(5)(450));
F6451: entity F port map(lamdaA => P(6)(451),lamdaB => P(6)(459),lamdaOut => P(5)(451));
F6452: entity F port map(lamdaA => P(6)(452),lamdaB => P(6)(460),lamdaOut => P(5)(452));
F6453: entity F port map(lamdaA => P(6)(453),lamdaB => P(6)(461),lamdaOut => P(5)(453));
F6454: entity F port map(lamdaA => P(6)(454),lamdaB => P(6)(462),lamdaOut => P(5)(454));
F6455: entity F port map(lamdaA => P(6)(455),lamdaB => P(6)(463),lamdaOut => P(5)(455));
G6456: entity G port map(lamdaA => P(6)(448),lamdaB => P(6)(456),s => s(6)(224),lamdaOut => P(5)(456));
G6457: entity G port map(lamdaA => P(6)(449),lamdaB => P(6)(457),s => s(6)(225),lamdaOut => P(5)(457));
G6458: entity G port map(lamdaA => P(6)(450),lamdaB => P(6)(458),s => s(6)(226),lamdaOut => P(5)(458));
G6459: entity G port map(lamdaA => P(6)(451),lamdaB => P(6)(459),s => s(6)(227),lamdaOut => P(5)(459));
G6460: entity G port map(lamdaA => P(6)(452),lamdaB => P(6)(460),s => s(6)(228),lamdaOut => P(5)(460));
G6461: entity G port map(lamdaA => P(6)(453),lamdaB => P(6)(461),s => s(6)(229),lamdaOut => P(5)(461));
G6462: entity G port map(lamdaA => P(6)(454),lamdaB => P(6)(462),s => s(6)(230),lamdaOut => P(5)(462));
G6463: entity G port map(lamdaA => P(6)(455),lamdaB => P(6)(463),s => s(6)(231),lamdaOut => P(5)(463));
F6464: entity F port map(lamdaA => P(6)(464),lamdaB => P(6)(472),lamdaOut => P(5)(464));
F6465: entity F port map(lamdaA => P(6)(465),lamdaB => P(6)(473),lamdaOut => P(5)(465));
F6466: entity F port map(lamdaA => P(6)(466),lamdaB => P(6)(474),lamdaOut => P(5)(466));
F6467: entity F port map(lamdaA => P(6)(467),lamdaB => P(6)(475),lamdaOut => P(5)(467));
F6468: entity F port map(lamdaA => P(6)(468),lamdaB => P(6)(476),lamdaOut => P(5)(468));
F6469: entity F port map(lamdaA => P(6)(469),lamdaB => P(6)(477),lamdaOut => P(5)(469));
F6470: entity F port map(lamdaA => P(6)(470),lamdaB => P(6)(478),lamdaOut => P(5)(470));
F6471: entity F port map(lamdaA => P(6)(471),lamdaB => P(6)(479),lamdaOut => P(5)(471));
G6472: entity G port map(lamdaA => P(6)(464),lamdaB => P(6)(472),s => s(6)(232),lamdaOut => P(5)(472));
G6473: entity G port map(lamdaA => P(6)(465),lamdaB => P(6)(473),s => s(6)(233),lamdaOut => P(5)(473));
G6474: entity G port map(lamdaA => P(6)(466),lamdaB => P(6)(474),s => s(6)(234),lamdaOut => P(5)(474));
G6475: entity G port map(lamdaA => P(6)(467),lamdaB => P(6)(475),s => s(6)(235),lamdaOut => P(5)(475));
G6476: entity G port map(lamdaA => P(6)(468),lamdaB => P(6)(476),s => s(6)(236),lamdaOut => P(5)(476));
G6477: entity G port map(lamdaA => P(6)(469),lamdaB => P(6)(477),s => s(6)(237),lamdaOut => P(5)(477));
G6478: entity G port map(lamdaA => P(6)(470),lamdaB => P(6)(478),s => s(6)(238),lamdaOut => P(5)(478));
G6479: entity G port map(lamdaA => P(6)(471),lamdaB => P(6)(479),s => s(6)(239),lamdaOut => P(5)(479));
F6480: entity F port map(lamdaA => P(6)(480),lamdaB => P(6)(488),lamdaOut => P(5)(480));
F6481: entity F port map(lamdaA => P(6)(481),lamdaB => P(6)(489),lamdaOut => P(5)(481));
F6482: entity F port map(lamdaA => P(6)(482),lamdaB => P(6)(490),lamdaOut => P(5)(482));
F6483: entity F port map(lamdaA => P(6)(483),lamdaB => P(6)(491),lamdaOut => P(5)(483));
F6484: entity F port map(lamdaA => P(6)(484),lamdaB => P(6)(492),lamdaOut => P(5)(484));
F6485: entity F port map(lamdaA => P(6)(485),lamdaB => P(6)(493),lamdaOut => P(5)(485));
F6486: entity F port map(lamdaA => P(6)(486),lamdaB => P(6)(494),lamdaOut => P(5)(486));
F6487: entity F port map(lamdaA => P(6)(487),lamdaB => P(6)(495),lamdaOut => P(5)(487));
G6488: entity G port map(lamdaA => P(6)(480),lamdaB => P(6)(488),s => s(6)(240),lamdaOut => P(5)(488));
G6489: entity G port map(lamdaA => P(6)(481),lamdaB => P(6)(489),s => s(6)(241),lamdaOut => P(5)(489));
G6490: entity G port map(lamdaA => P(6)(482),lamdaB => P(6)(490),s => s(6)(242),lamdaOut => P(5)(490));
G6491: entity G port map(lamdaA => P(6)(483),lamdaB => P(6)(491),s => s(6)(243),lamdaOut => P(5)(491));
G6492: entity G port map(lamdaA => P(6)(484),lamdaB => P(6)(492),s => s(6)(244),lamdaOut => P(5)(492));
G6493: entity G port map(lamdaA => P(6)(485),lamdaB => P(6)(493),s => s(6)(245),lamdaOut => P(5)(493));
G6494: entity G port map(lamdaA => P(6)(486),lamdaB => P(6)(494),s => s(6)(246),lamdaOut => P(5)(494));
G6495: entity G port map(lamdaA => P(6)(487),lamdaB => P(6)(495),s => s(6)(247),lamdaOut => P(5)(495));
F6496: entity F port map(lamdaA => P(6)(496),lamdaB => P(6)(504),lamdaOut => P(5)(496));
F6497: entity F port map(lamdaA => P(6)(497),lamdaB => P(6)(505),lamdaOut => P(5)(497));
F6498: entity F port map(lamdaA => P(6)(498),lamdaB => P(6)(506),lamdaOut => P(5)(498));
F6499: entity F port map(lamdaA => P(6)(499),lamdaB => P(6)(507),lamdaOut => P(5)(499));
F6500: entity F port map(lamdaA => P(6)(500),lamdaB => P(6)(508),lamdaOut => P(5)(500));
F6501: entity F port map(lamdaA => P(6)(501),lamdaB => P(6)(509),lamdaOut => P(5)(501));
F6502: entity F port map(lamdaA => P(6)(502),lamdaB => P(6)(510),lamdaOut => P(5)(502));
F6503: entity F port map(lamdaA => P(6)(503),lamdaB => P(6)(511),lamdaOut => P(5)(503));
G6504: entity G port map(lamdaA => P(6)(496),lamdaB => P(6)(504),s => s(6)(248),lamdaOut => P(5)(504));
G6505: entity G port map(lamdaA => P(6)(497),lamdaB => P(6)(505),s => s(6)(249),lamdaOut => P(5)(505));
G6506: entity G port map(lamdaA => P(6)(498),lamdaB => P(6)(506),s => s(6)(250),lamdaOut => P(5)(506));
G6507: entity G port map(lamdaA => P(6)(499),lamdaB => P(6)(507),s => s(6)(251),lamdaOut => P(5)(507));
G6508: entity G port map(lamdaA => P(6)(500),lamdaB => P(6)(508),s => s(6)(252),lamdaOut => P(5)(508));
G6509: entity G port map(lamdaA => P(6)(501),lamdaB => P(6)(509),s => s(6)(253),lamdaOut => P(5)(509));
G6510: entity G port map(lamdaA => P(6)(502),lamdaB => P(6)(510),s => s(6)(254),lamdaOut => P(5)(510));
G6511: entity G port map(lamdaA => P(6)(503),lamdaB => P(6)(511),s => s(6)(255),lamdaOut => P(5)(511));
-- STAGE 5
F50: entity F port map(lamdaA => P(5)(0),lamdaB => P(5)(16),lamdaOut => P(4)(0));
F51: entity F port map(lamdaA => P(5)(1),lamdaB => P(5)(17),lamdaOut => P(4)(1));
F52: entity F port map(lamdaA => P(5)(2),lamdaB => P(5)(18),lamdaOut => P(4)(2));
F53: entity F port map(lamdaA => P(5)(3),lamdaB => P(5)(19),lamdaOut => P(4)(3));
F54: entity F port map(lamdaA => P(5)(4),lamdaB => P(5)(20),lamdaOut => P(4)(4));
F55: entity F port map(lamdaA => P(5)(5),lamdaB => P(5)(21),lamdaOut => P(4)(5));
F56: entity F port map(lamdaA => P(5)(6),lamdaB => P(5)(22),lamdaOut => P(4)(6));
F57: entity F port map(lamdaA => P(5)(7),lamdaB => P(5)(23),lamdaOut => P(4)(7));
F58: entity F port map(lamdaA => P(5)(8),lamdaB => P(5)(24),lamdaOut => P(4)(8));
F59: entity F port map(lamdaA => P(5)(9),lamdaB => P(5)(25),lamdaOut => P(4)(9));
F510: entity F port map(lamdaA => P(5)(10),lamdaB => P(5)(26),lamdaOut => P(4)(10));
F511: entity F port map(lamdaA => P(5)(11),lamdaB => P(5)(27),lamdaOut => P(4)(11));
F512: entity F port map(lamdaA => P(5)(12),lamdaB => P(5)(28),lamdaOut => P(4)(12));
F513: entity F port map(lamdaA => P(5)(13),lamdaB => P(5)(29),lamdaOut => P(4)(13));
F514: entity F port map(lamdaA => P(5)(14),lamdaB => P(5)(30),lamdaOut => P(4)(14));
F515: entity F port map(lamdaA => P(5)(15),lamdaB => P(5)(31),lamdaOut => P(4)(15));
G516: entity G port map(lamdaA => P(5)(0),lamdaB => P(5)(16),s => s(5)(0),lamdaOut => P(4)(16));
G517: entity G port map(lamdaA => P(5)(1),lamdaB => P(5)(17),s => s(5)(1),lamdaOut => P(4)(17));
G518: entity G port map(lamdaA => P(5)(2),lamdaB => P(5)(18),s => s(5)(2),lamdaOut => P(4)(18));
G519: entity G port map(lamdaA => P(5)(3),lamdaB => P(5)(19),s => s(5)(3),lamdaOut => P(4)(19));
G520: entity G port map(lamdaA => P(5)(4),lamdaB => P(5)(20),s => s(5)(4),lamdaOut => P(4)(20));
G521: entity G port map(lamdaA => P(5)(5),lamdaB => P(5)(21),s => s(5)(5),lamdaOut => P(4)(21));
G522: entity G port map(lamdaA => P(5)(6),lamdaB => P(5)(22),s => s(5)(6),lamdaOut => P(4)(22));
G523: entity G port map(lamdaA => P(5)(7),lamdaB => P(5)(23),s => s(5)(7),lamdaOut => P(4)(23));
G524: entity G port map(lamdaA => P(5)(8),lamdaB => P(5)(24),s => s(5)(8),lamdaOut => P(4)(24));
G525: entity G port map(lamdaA => P(5)(9),lamdaB => P(5)(25),s => s(5)(9),lamdaOut => P(4)(25));
G526: entity G port map(lamdaA => P(5)(10),lamdaB => P(5)(26),s => s(5)(10),lamdaOut => P(4)(26));
G527: entity G port map(lamdaA => P(5)(11),lamdaB => P(5)(27),s => s(5)(11),lamdaOut => P(4)(27));
G528: entity G port map(lamdaA => P(5)(12),lamdaB => P(5)(28),s => s(5)(12),lamdaOut => P(4)(28));
G529: entity G port map(lamdaA => P(5)(13),lamdaB => P(5)(29),s => s(5)(13),lamdaOut => P(4)(29));
G530: entity G port map(lamdaA => P(5)(14),lamdaB => P(5)(30),s => s(5)(14),lamdaOut => P(4)(30));
G531: entity G port map(lamdaA => P(5)(15),lamdaB => P(5)(31),s => s(5)(15),lamdaOut => P(4)(31));
F532: entity F port map(lamdaA => P(5)(32),lamdaB => P(5)(48),lamdaOut => P(4)(32));
F533: entity F port map(lamdaA => P(5)(33),lamdaB => P(5)(49),lamdaOut => P(4)(33));
F534: entity F port map(lamdaA => P(5)(34),lamdaB => P(5)(50),lamdaOut => P(4)(34));
F535: entity F port map(lamdaA => P(5)(35),lamdaB => P(5)(51),lamdaOut => P(4)(35));
F536: entity F port map(lamdaA => P(5)(36),lamdaB => P(5)(52),lamdaOut => P(4)(36));
F537: entity F port map(lamdaA => P(5)(37),lamdaB => P(5)(53),lamdaOut => P(4)(37));
F538: entity F port map(lamdaA => P(5)(38),lamdaB => P(5)(54),lamdaOut => P(4)(38));
F539: entity F port map(lamdaA => P(5)(39),lamdaB => P(5)(55),lamdaOut => P(4)(39));
F540: entity F port map(lamdaA => P(5)(40),lamdaB => P(5)(56),lamdaOut => P(4)(40));
F541: entity F port map(lamdaA => P(5)(41),lamdaB => P(5)(57),lamdaOut => P(4)(41));
F542: entity F port map(lamdaA => P(5)(42),lamdaB => P(5)(58),lamdaOut => P(4)(42));
F543: entity F port map(lamdaA => P(5)(43),lamdaB => P(5)(59),lamdaOut => P(4)(43));
F544: entity F port map(lamdaA => P(5)(44),lamdaB => P(5)(60),lamdaOut => P(4)(44));
F545: entity F port map(lamdaA => P(5)(45),lamdaB => P(5)(61),lamdaOut => P(4)(45));
F546: entity F port map(lamdaA => P(5)(46),lamdaB => P(5)(62),lamdaOut => P(4)(46));
F547: entity F port map(lamdaA => P(5)(47),lamdaB => P(5)(63),lamdaOut => P(4)(47));
G548: entity G port map(lamdaA => P(5)(32),lamdaB => P(5)(48),s => s(5)(16),lamdaOut => P(4)(48));
G549: entity G port map(lamdaA => P(5)(33),lamdaB => P(5)(49),s => s(5)(17),lamdaOut => P(4)(49));
G550: entity G port map(lamdaA => P(5)(34),lamdaB => P(5)(50),s => s(5)(18),lamdaOut => P(4)(50));
G551: entity G port map(lamdaA => P(5)(35),lamdaB => P(5)(51),s => s(5)(19),lamdaOut => P(4)(51));
G552: entity G port map(lamdaA => P(5)(36),lamdaB => P(5)(52),s => s(5)(20),lamdaOut => P(4)(52));
G553: entity G port map(lamdaA => P(5)(37),lamdaB => P(5)(53),s => s(5)(21),lamdaOut => P(4)(53));
G554: entity G port map(lamdaA => P(5)(38),lamdaB => P(5)(54),s => s(5)(22),lamdaOut => P(4)(54));
G555: entity G port map(lamdaA => P(5)(39),lamdaB => P(5)(55),s => s(5)(23),lamdaOut => P(4)(55));
G556: entity G port map(lamdaA => P(5)(40),lamdaB => P(5)(56),s => s(5)(24),lamdaOut => P(4)(56));
G557: entity G port map(lamdaA => P(5)(41),lamdaB => P(5)(57),s => s(5)(25),lamdaOut => P(4)(57));
G558: entity G port map(lamdaA => P(5)(42),lamdaB => P(5)(58),s => s(5)(26),lamdaOut => P(4)(58));
G559: entity G port map(lamdaA => P(5)(43),lamdaB => P(5)(59),s => s(5)(27),lamdaOut => P(4)(59));
G560: entity G port map(lamdaA => P(5)(44),lamdaB => P(5)(60),s => s(5)(28),lamdaOut => P(4)(60));
G561: entity G port map(lamdaA => P(5)(45),lamdaB => P(5)(61),s => s(5)(29),lamdaOut => P(4)(61));
G562: entity G port map(lamdaA => P(5)(46),lamdaB => P(5)(62),s => s(5)(30),lamdaOut => P(4)(62));
G563: entity G port map(lamdaA => P(5)(47),lamdaB => P(5)(63),s => s(5)(31),lamdaOut => P(4)(63));
F564: entity F port map(lamdaA => P(5)(64),lamdaB => P(5)(80),lamdaOut => P(4)(64));
F565: entity F port map(lamdaA => P(5)(65),lamdaB => P(5)(81),lamdaOut => P(4)(65));
F566: entity F port map(lamdaA => P(5)(66),lamdaB => P(5)(82),lamdaOut => P(4)(66));
F567: entity F port map(lamdaA => P(5)(67),lamdaB => P(5)(83),lamdaOut => P(4)(67));
F568: entity F port map(lamdaA => P(5)(68),lamdaB => P(5)(84),lamdaOut => P(4)(68));
F569: entity F port map(lamdaA => P(5)(69),lamdaB => P(5)(85),lamdaOut => P(4)(69));
F570: entity F port map(lamdaA => P(5)(70),lamdaB => P(5)(86),lamdaOut => P(4)(70));
F571: entity F port map(lamdaA => P(5)(71),lamdaB => P(5)(87),lamdaOut => P(4)(71));
F572: entity F port map(lamdaA => P(5)(72),lamdaB => P(5)(88),lamdaOut => P(4)(72));
F573: entity F port map(lamdaA => P(5)(73),lamdaB => P(5)(89),lamdaOut => P(4)(73));
F574: entity F port map(lamdaA => P(5)(74),lamdaB => P(5)(90),lamdaOut => P(4)(74));
F575: entity F port map(lamdaA => P(5)(75),lamdaB => P(5)(91),lamdaOut => P(4)(75));
F576: entity F port map(lamdaA => P(5)(76),lamdaB => P(5)(92),lamdaOut => P(4)(76));
F577: entity F port map(lamdaA => P(5)(77),lamdaB => P(5)(93),lamdaOut => P(4)(77));
F578: entity F port map(lamdaA => P(5)(78),lamdaB => P(5)(94),lamdaOut => P(4)(78));
F579: entity F port map(lamdaA => P(5)(79),lamdaB => P(5)(95),lamdaOut => P(4)(79));
G580: entity G port map(lamdaA => P(5)(64),lamdaB => P(5)(80),s => s(5)(32),lamdaOut => P(4)(80));
G581: entity G port map(lamdaA => P(5)(65),lamdaB => P(5)(81),s => s(5)(33),lamdaOut => P(4)(81));
G582: entity G port map(lamdaA => P(5)(66),lamdaB => P(5)(82),s => s(5)(34),lamdaOut => P(4)(82));
G583: entity G port map(lamdaA => P(5)(67),lamdaB => P(5)(83),s => s(5)(35),lamdaOut => P(4)(83));
G584: entity G port map(lamdaA => P(5)(68),lamdaB => P(5)(84),s => s(5)(36),lamdaOut => P(4)(84));
G585: entity G port map(lamdaA => P(5)(69),lamdaB => P(5)(85),s => s(5)(37),lamdaOut => P(4)(85));
G586: entity G port map(lamdaA => P(5)(70),lamdaB => P(5)(86),s => s(5)(38),lamdaOut => P(4)(86));
G587: entity G port map(lamdaA => P(5)(71),lamdaB => P(5)(87),s => s(5)(39),lamdaOut => P(4)(87));
G588: entity G port map(lamdaA => P(5)(72),lamdaB => P(5)(88),s => s(5)(40),lamdaOut => P(4)(88));
G589: entity G port map(lamdaA => P(5)(73),lamdaB => P(5)(89),s => s(5)(41),lamdaOut => P(4)(89));
G590: entity G port map(lamdaA => P(5)(74),lamdaB => P(5)(90),s => s(5)(42),lamdaOut => P(4)(90));
G591: entity G port map(lamdaA => P(5)(75),lamdaB => P(5)(91),s => s(5)(43),lamdaOut => P(4)(91));
G592: entity G port map(lamdaA => P(5)(76),lamdaB => P(5)(92),s => s(5)(44),lamdaOut => P(4)(92));
G593: entity G port map(lamdaA => P(5)(77),lamdaB => P(5)(93),s => s(5)(45),lamdaOut => P(4)(93));
G594: entity G port map(lamdaA => P(5)(78),lamdaB => P(5)(94),s => s(5)(46),lamdaOut => P(4)(94));
G595: entity G port map(lamdaA => P(5)(79),lamdaB => P(5)(95),s => s(5)(47),lamdaOut => P(4)(95));
F596: entity F port map(lamdaA => P(5)(96),lamdaB => P(5)(112),lamdaOut => P(4)(96));
F597: entity F port map(lamdaA => P(5)(97),lamdaB => P(5)(113),lamdaOut => P(4)(97));
F598: entity F port map(lamdaA => P(5)(98),lamdaB => P(5)(114),lamdaOut => P(4)(98));
F599: entity F port map(lamdaA => P(5)(99),lamdaB => P(5)(115),lamdaOut => P(4)(99));
F5100: entity F port map(lamdaA => P(5)(100),lamdaB => P(5)(116),lamdaOut => P(4)(100));
F5101: entity F port map(lamdaA => P(5)(101),lamdaB => P(5)(117),lamdaOut => P(4)(101));
F5102: entity F port map(lamdaA => P(5)(102),lamdaB => P(5)(118),lamdaOut => P(4)(102));
F5103: entity F port map(lamdaA => P(5)(103),lamdaB => P(5)(119),lamdaOut => P(4)(103));
F5104: entity F port map(lamdaA => P(5)(104),lamdaB => P(5)(120),lamdaOut => P(4)(104));
F5105: entity F port map(lamdaA => P(5)(105),lamdaB => P(5)(121),lamdaOut => P(4)(105));
F5106: entity F port map(lamdaA => P(5)(106),lamdaB => P(5)(122),lamdaOut => P(4)(106));
F5107: entity F port map(lamdaA => P(5)(107),lamdaB => P(5)(123),lamdaOut => P(4)(107));
F5108: entity F port map(lamdaA => P(5)(108),lamdaB => P(5)(124),lamdaOut => P(4)(108));
F5109: entity F port map(lamdaA => P(5)(109),lamdaB => P(5)(125),lamdaOut => P(4)(109));
F5110: entity F port map(lamdaA => P(5)(110),lamdaB => P(5)(126),lamdaOut => P(4)(110));
F5111: entity F port map(lamdaA => P(5)(111),lamdaB => P(5)(127),lamdaOut => P(4)(111));
G5112: entity G port map(lamdaA => P(5)(96),lamdaB => P(5)(112),s => s(5)(48),lamdaOut => P(4)(112));
G5113: entity G port map(lamdaA => P(5)(97),lamdaB => P(5)(113),s => s(5)(49),lamdaOut => P(4)(113));
G5114: entity G port map(lamdaA => P(5)(98),lamdaB => P(5)(114),s => s(5)(50),lamdaOut => P(4)(114));
G5115: entity G port map(lamdaA => P(5)(99),lamdaB => P(5)(115),s => s(5)(51),lamdaOut => P(4)(115));
G5116: entity G port map(lamdaA => P(5)(100),lamdaB => P(5)(116),s => s(5)(52),lamdaOut => P(4)(116));
G5117: entity G port map(lamdaA => P(5)(101),lamdaB => P(5)(117),s => s(5)(53),lamdaOut => P(4)(117));
G5118: entity G port map(lamdaA => P(5)(102),lamdaB => P(5)(118),s => s(5)(54),lamdaOut => P(4)(118));
G5119: entity G port map(lamdaA => P(5)(103),lamdaB => P(5)(119),s => s(5)(55),lamdaOut => P(4)(119));
G5120: entity G port map(lamdaA => P(5)(104),lamdaB => P(5)(120),s => s(5)(56),lamdaOut => P(4)(120));
G5121: entity G port map(lamdaA => P(5)(105),lamdaB => P(5)(121),s => s(5)(57),lamdaOut => P(4)(121));
G5122: entity G port map(lamdaA => P(5)(106),lamdaB => P(5)(122),s => s(5)(58),lamdaOut => P(4)(122));
G5123: entity G port map(lamdaA => P(5)(107),lamdaB => P(5)(123),s => s(5)(59),lamdaOut => P(4)(123));
G5124: entity G port map(lamdaA => P(5)(108),lamdaB => P(5)(124),s => s(5)(60),lamdaOut => P(4)(124));
G5125: entity G port map(lamdaA => P(5)(109),lamdaB => P(5)(125),s => s(5)(61),lamdaOut => P(4)(125));
G5126: entity G port map(lamdaA => P(5)(110),lamdaB => P(5)(126),s => s(5)(62),lamdaOut => P(4)(126));
G5127: entity G port map(lamdaA => P(5)(111),lamdaB => P(5)(127),s => s(5)(63),lamdaOut => P(4)(127));
F5128: entity F port map(lamdaA => P(5)(128),lamdaB => P(5)(144),lamdaOut => P(4)(128));
F5129: entity F port map(lamdaA => P(5)(129),lamdaB => P(5)(145),lamdaOut => P(4)(129));
F5130: entity F port map(lamdaA => P(5)(130),lamdaB => P(5)(146),lamdaOut => P(4)(130));
F5131: entity F port map(lamdaA => P(5)(131),lamdaB => P(5)(147),lamdaOut => P(4)(131));
F5132: entity F port map(lamdaA => P(5)(132),lamdaB => P(5)(148),lamdaOut => P(4)(132));
F5133: entity F port map(lamdaA => P(5)(133),lamdaB => P(5)(149),lamdaOut => P(4)(133));
F5134: entity F port map(lamdaA => P(5)(134),lamdaB => P(5)(150),lamdaOut => P(4)(134));
F5135: entity F port map(lamdaA => P(5)(135),lamdaB => P(5)(151),lamdaOut => P(4)(135));
F5136: entity F port map(lamdaA => P(5)(136),lamdaB => P(5)(152),lamdaOut => P(4)(136));
F5137: entity F port map(lamdaA => P(5)(137),lamdaB => P(5)(153),lamdaOut => P(4)(137));
F5138: entity F port map(lamdaA => P(5)(138),lamdaB => P(5)(154),lamdaOut => P(4)(138));
F5139: entity F port map(lamdaA => P(5)(139),lamdaB => P(5)(155),lamdaOut => P(4)(139));
F5140: entity F port map(lamdaA => P(5)(140),lamdaB => P(5)(156),lamdaOut => P(4)(140));
F5141: entity F port map(lamdaA => P(5)(141),lamdaB => P(5)(157),lamdaOut => P(4)(141));
F5142: entity F port map(lamdaA => P(5)(142),lamdaB => P(5)(158),lamdaOut => P(4)(142));
F5143: entity F port map(lamdaA => P(5)(143),lamdaB => P(5)(159),lamdaOut => P(4)(143));
G5144: entity G port map(lamdaA => P(5)(128),lamdaB => P(5)(144),s => s(5)(64),lamdaOut => P(4)(144));
G5145: entity G port map(lamdaA => P(5)(129),lamdaB => P(5)(145),s => s(5)(65),lamdaOut => P(4)(145));
G5146: entity G port map(lamdaA => P(5)(130),lamdaB => P(5)(146),s => s(5)(66),lamdaOut => P(4)(146));
G5147: entity G port map(lamdaA => P(5)(131),lamdaB => P(5)(147),s => s(5)(67),lamdaOut => P(4)(147));
G5148: entity G port map(lamdaA => P(5)(132),lamdaB => P(5)(148),s => s(5)(68),lamdaOut => P(4)(148));
G5149: entity G port map(lamdaA => P(5)(133),lamdaB => P(5)(149),s => s(5)(69),lamdaOut => P(4)(149));
G5150: entity G port map(lamdaA => P(5)(134),lamdaB => P(5)(150),s => s(5)(70),lamdaOut => P(4)(150));
G5151: entity G port map(lamdaA => P(5)(135),lamdaB => P(5)(151),s => s(5)(71),lamdaOut => P(4)(151));
G5152: entity G port map(lamdaA => P(5)(136),lamdaB => P(5)(152),s => s(5)(72),lamdaOut => P(4)(152));
G5153: entity G port map(lamdaA => P(5)(137),lamdaB => P(5)(153),s => s(5)(73),lamdaOut => P(4)(153));
G5154: entity G port map(lamdaA => P(5)(138),lamdaB => P(5)(154),s => s(5)(74),lamdaOut => P(4)(154));
G5155: entity G port map(lamdaA => P(5)(139),lamdaB => P(5)(155),s => s(5)(75),lamdaOut => P(4)(155));
G5156: entity G port map(lamdaA => P(5)(140),lamdaB => P(5)(156),s => s(5)(76),lamdaOut => P(4)(156));
G5157: entity G port map(lamdaA => P(5)(141),lamdaB => P(5)(157),s => s(5)(77),lamdaOut => P(4)(157));
G5158: entity G port map(lamdaA => P(5)(142),lamdaB => P(5)(158),s => s(5)(78),lamdaOut => P(4)(158));
G5159: entity G port map(lamdaA => P(5)(143),lamdaB => P(5)(159),s => s(5)(79),lamdaOut => P(4)(159));
F5160: entity F port map(lamdaA => P(5)(160),lamdaB => P(5)(176),lamdaOut => P(4)(160));
F5161: entity F port map(lamdaA => P(5)(161),lamdaB => P(5)(177),lamdaOut => P(4)(161));
F5162: entity F port map(lamdaA => P(5)(162),lamdaB => P(5)(178),lamdaOut => P(4)(162));
F5163: entity F port map(lamdaA => P(5)(163),lamdaB => P(5)(179),lamdaOut => P(4)(163));
F5164: entity F port map(lamdaA => P(5)(164),lamdaB => P(5)(180),lamdaOut => P(4)(164));
F5165: entity F port map(lamdaA => P(5)(165),lamdaB => P(5)(181),lamdaOut => P(4)(165));
F5166: entity F port map(lamdaA => P(5)(166),lamdaB => P(5)(182),lamdaOut => P(4)(166));
F5167: entity F port map(lamdaA => P(5)(167),lamdaB => P(5)(183),lamdaOut => P(4)(167));
F5168: entity F port map(lamdaA => P(5)(168),lamdaB => P(5)(184),lamdaOut => P(4)(168));
F5169: entity F port map(lamdaA => P(5)(169),lamdaB => P(5)(185),lamdaOut => P(4)(169));
F5170: entity F port map(lamdaA => P(5)(170),lamdaB => P(5)(186),lamdaOut => P(4)(170));
F5171: entity F port map(lamdaA => P(5)(171),lamdaB => P(5)(187),lamdaOut => P(4)(171));
F5172: entity F port map(lamdaA => P(5)(172),lamdaB => P(5)(188),lamdaOut => P(4)(172));
F5173: entity F port map(lamdaA => P(5)(173),lamdaB => P(5)(189),lamdaOut => P(4)(173));
F5174: entity F port map(lamdaA => P(5)(174),lamdaB => P(5)(190),lamdaOut => P(4)(174));
F5175: entity F port map(lamdaA => P(5)(175),lamdaB => P(5)(191),lamdaOut => P(4)(175));
G5176: entity G port map(lamdaA => P(5)(160),lamdaB => P(5)(176),s => s(5)(80),lamdaOut => P(4)(176));
G5177: entity G port map(lamdaA => P(5)(161),lamdaB => P(5)(177),s => s(5)(81),lamdaOut => P(4)(177));
G5178: entity G port map(lamdaA => P(5)(162),lamdaB => P(5)(178),s => s(5)(82),lamdaOut => P(4)(178));
G5179: entity G port map(lamdaA => P(5)(163),lamdaB => P(5)(179),s => s(5)(83),lamdaOut => P(4)(179));
G5180: entity G port map(lamdaA => P(5)(164),lamdaB => P(5)(180),s => s(5)(84),lamdaOut => P(4)(180));
G5181: entity G port map(lamdaA => P(5)(165),lamdaB => P(5)(181),s => s(5)(85),lamdaOut => P(4)(181));
G5182: entity G port map(lamdaA => P(5)(166),lamdaB => P(5)(182),s => s(5)(86),lamdaOut => P(4)(182));
G5183: entity G port map(lamdaA => P(5)(167),lamdaB => P(5)(183),s => s(5)(87),lamdaOut => P(4)(183));
G5184: entity G port map(lamdaA => P(5)(168),lamdaB => P(5)(184),s => s(5)(88),lamdaOut => P(4)(184));
G5185: entity G port map(lamdaA => P(5)(169),lamdaB => P(5)(185),s => s(5)(89),lamdaOut => P(4)(185));
G5186: entity G port map(lamdaA => P(5)(170),lamdaB => P(5)(186),s => s(5)(90),lamdaOut => P(4)(186));
G5187: entity G port map(lamdaA => P(5)(171),lamdaB => P(5)(187),s => s(5)(91),lamdaOut => P(4)(187));
G5188: entity G port map(lamdaA => P(5)(172),lamdaB => P(5)(188),s => s(5)(92),lamdaOut => P(4)(188));
G5189: entity G port map(lamdaA => P(5)(173),lamdaB => P(5)(189),s => s(5)(93),lamdaOut => P(4)(189));
G5190: entity G port map(lamdaA => P(5)(174),lamdaB => P(5)(190),s => s(5)(94),lamdaOut => P(4)(190));
G5191: entity G port map(lamdaA => P(5)(175),lamdaB => P(5)(191),s => s(5)(95),lamdaOut => P(4)(191));
F5192: entity F port map(lamdaA => P(5)(192),lamdaB => P(5)(208),lamdaOut => P(4)(192));
F5193: entity F port map(lamdaA => P(5)(193),lamdaB => P(5)(209),lamdaOut => P(4)(193));
F5194: entity F port map(lamdaA => P(5)(194),lamdaB => P(5)(210),lamdaOut => P(4)(194));
F5195: entity F port map(lamdaA => P(5)(195),lamdaB => P(5)(211),lamdaOut => P(4)(195));
F5196: entity F port map(lamdaA => P(5)(196),lamdaB => P(5)(212),lamdaOut => P(4)(196));
F5197: entity F port map(lamdaA => P(5)(197),lamdaB => P(5)(213),lamdaOut => P(4)(197));
F5198: entity F port map(lamdaA => P(5)(198),lamdaB => P(5)(214),lamdaOut => P(4)(198));
F5199: entity F port map(lamdaA => P(5)(199),lamdaB => P(5)(215),lamdaOut => P(4)(199));
F5200: entity F port map(lamdaA => P(5)(200),lamdaB => P(5)(216),lamdaOut => P(4)(200));
F5201: entity F port map(lamdaA => P(5)(201),lamdaB => P(5)(217),lamdaOut => P(4)(201));
F5202: entity F port map(lamdaA => P(5)(202),lamdaB => P(5)(218),lamdaOut => P(4)(202));
F5203: entity F port map(lamdaA => P(5)(203),lamdaB => P(5)(219),lamdaOut => P(4)(203));
F5204: entity F port map(lamdaA => P(5)(204),lamdaB => P(5)(220),lamdaOut => P(4)(204));
F5205: entity F port map(lamdaA => P(5)(205),lamdaB => P(5)(221),lamdaOut => P(4)(205));
F5206: entity F port map(lamdaA => P(5)(206),lamdaB => P(5)(222),lamdaOut => P(4)(206));
F5207: entity F port map(lamdaA => P(5)(207),lamdaB => P(5)(223),lamdaOut => P(4)(207));
G5208: entity G port map(lamdaA => P(5)(192),lamdaB => P(5)(208),s => s(5)(96),lamdaOut => P(4)(208));
G5209: entity G port map(lamdaA => P(5)(193),lamdaB => P(5)(209),s => s(5)(97),lamdaOut => P(4)(209));
G5210: entity G port map(lamdaA => P(5)(194),lamdaB => P(5)(210),s => s(5)(98),lamdaOut => P(4)(210));
G5211: entity G port map(lamdaA => P(5)(195),lamdaB => P(5)(211),s => s(5)(99),lamdaOut => P(4)(211));
G5212: entity G port map(lamdaA => P(5)(196),lamdaB => P(5)(212),s => s(5)(100),lamdaOut => P(4)(212));
G5213: entity G port map(lamdaA => P(5)(197),lamdaB => P(5)(213),s => s(5)(101),lamdaOut => P(4)(213));
G5214: entity G port map(lamdaA => P(5)(198),lamdaB => P(5)(214),s => s(5)(102),lamdaOut => P(4)(214));
G5215: entity G port map(lamdaA => P(5)(199),lamdaB => P(5)(215),s => s(5)(103),lamdaOut => P(4)(215));
G5216: entity G port map(lamdaA => P(5)(200),lamdaB => P(5)(216),s => s(5)(104),lamdaOut => P(4)(216));
G5217: entity G port map(lamdaA => P(5)(201),lamdaB => P(5)(217),s => s(5)(105),lamdaOut => P(4)(217));
G5218: entity G port map(lamdaA => P(5)(202),lamdaB => P(5)(218),s => s(5)(106),lamdaOut => P(4)(218));
G5219: entity G port map(lamdaA => P(5)(203),lamdaB => P(5)(219),s => s(5)(107),lamdaOut => P(4)(219));
G5220: entity G port map(lamdaA => P(5)(204),lamdaB => P(5)(220),s => s(5)(108),lamdaOut => P(4)(220));
G5221: entity G port map(lamdaA => P(5)(205),lamdaB => P(5)(221),s => s(5)(109),lamdaOut => P(4)(221));
G5222: entity G port map(lamdaA => P(5)(206),lamdaB => P(5)(222),s => s(5)(110),lamdaOut => P(4)(222));
G5223: entity G port map(lamdaA => P(5)(207),lamdaB => P(5)(223),s => s(5)(111),lamdaOut => P(4)(223));
F5224: entity F port map(lamdaA => P(5)(224),lamdaB => P(5)(240),lamdaOut => P(4)(224));
F5225: entity F port map(lamdaA => P(5)(225),lamdaB => P(5)(241),lamdaOut => P(4)(225));
F5226: entity F port map(lamdaA => P(5)(226),lamdaB => P(5)(242),lamdaOut => P(4)(226));
F5227: entity F port map(lamdaA => P(5)(227),lamdaB => P(5)(243),lamdaOut => P(4)(227));
F5228: entity F port map(lamdaA => P(5)(228),lamdaB => P(5)(244),lamdaOut => P(4)(228));
F5229: entity F port map(lamdaA => P(5)(229),lamdaB => P(5)(245),lamdaOut => P(4)(229));
F5230: entity F port map(lamdaA => P(5)(230),lamdaB => P(5)(246),lamdaOut => P(4)(230));
F5231: entity F port map(lamdaA => P(5)(231),lamdaB => P(5)(247),lamdaOut => P(4)(231));
F5232: entity F port map(lamdaA => P(5)(232),lamdaB => P(5)(248),lamdaOut => P(4)(232));
F5233: entity F port map(lamdaA => P(5)(233),lamdaB => P(5)(249),lamdaOut => P(4)(233));
F5234: entity F port map(lamdaA => P(5)(234),lamdaB => P(5)(250),lamdaOut => P(4)(234));
F5235: entity F port map(lamdaA => P(5)(235),lamdaB => P(5)(251),lamdaOut => P(4)(235));
F5236: entity F port map(lamdaA => P(5)(236),lamdaB => P(5)(252),lamdaOut => P(4)(236));
F5237: entity F port map(lamdaA => P(5)(237),lamdaB => P(5)(253),lamdaOut => P(4)(237));
F5238: entity F port map(lamdaA => P(5)(238),lamdaB => P(5)(254),lamdaOut => P(4)(238));
F5239: entity F port map(lamdaA => P(5)(239),lamdaB => P(5)(255),lamdaOut => P(4)(239));
G5240: entity G port map(lamdaA => P(5)(224),lamdaB => P(5)(240),s => s(5)(112),lamdaOut => P(4)(240));
G5241: entity G port map(lamdaA => P(5)(225),lamdaB => P(5)(241),s => s(5)(113),lamdaOut => P(4)(241));
G5242: entity G port map(lamdaA => P(5)(226),lamdaB => P(5)(242),s => s(5)(114),lamdaOut => P(4)(242));
G5243: entity G port map(lamdaA => P(5)(227),lamdaB => P(5)(243),s => s(5)(115),lamdaOut => P(4)(243));
G5244: entity G port map(lamdaA => P(5)(228),lamdaB => P(5)(244),s => s(5)(116),lamdaOut => P(4)(244));
G5245: entity G port map(lamdaA => P(5)(229),lamdaB => P(5)(245),s => s(5)(117),lamdaOut => P(4)(245));
G5246: entity G port map(lamdaA => P(5)(230),lamdaB => P(5)(246),s => s(5)(118),lamdaOut => P(4)(246));
G5247: entity G port map(lamdaA => P(5)(231),lamdaB => P(5)(247),s => s(5)(119),lamdaOut => P(4)(247));
G5248: entity G port map(lamdaA => P(5)(232),lamdaB => P(5)(248),s => s(5)(120),lamdaOut => P(4)(248));
G5249: entity G port map(lamdaA => P(5)(233),lamdaB => P(5)(249),s => s(5)(121),lamdaOut => P(4)(249));
G5250: entity G port map(lamdaA => P(5)(234),lamdaB => P(5)(250),s => s(5)(122),lamdaOut => P(4)(250));
G5251: entity G port map(lamdaA => P(5)(235),lamdaB => P(5)(251),s => s(5)(123),lamdaOut => P(4)(251));
G5252: entity G port map(lamdaA => P(5)(236),lamdaB => P(5)(252),s => s(5)(124),lamdaOut => P(4)(252));
G5253: entity G port map(lamdaA => P(5)(237),lamdaB => P(5)(253),s => s(5)(125),lamdaOut => P(4)(253));
G5254: entity G port map(lamdaA => P(5)(238),lamdaB => P(5)(254),s => s(5)(126),lamdaOut => P(4)(254));
G5255: entity G port map(lamdaA => P(5)(239),lamdaB => P(5)(255),s => s(5)(127),lamdaOut => P(4)(255));
F5256: entity F port map(lamdaA => P(5)(256),lamdaB => P(5)(272),lamdaOut => P(4)(256));
F5257: entity F port map(lamdaA => P(5)(257),lamdaB => P(5)(273),lamdaOut => P(4)(257));
F5258: entity F port map(lamdaA => P(5)(258),lamdaB => P(5)(274),lamdaOut => P(4)(258));
F5259: entity F port map(lamdaA => P(5)(259),lamdaB => P(5)(275),lamdaOut => P(4)(259));
F5260: entity F port map(lamdaA => P(5)(260),lamdaB => P(5)(276),lamdaOut => P(4)(260));
F5261: entity F port map(lamdaA => P(5)(261),lamdaB => P(5)(277),lamdaOut => P(4)(261));
F5262: entity F port map(lamdaA => P(5)(262),lamdaB => P(5)(278),lamdaOut => P(4)(262));
F5263: entity F port map(lamdaA => P(5)(263),lamdaB => P(5)(279),lamdaOut => P(4)(263));
F5264: entity F port map(lamdaA => P(5)(264),lamdaB => P(5)(280),lamdaOut => P(4)(264));
F5265: entity F port map(lamdaA => P(5)(265),lamdaB => P(5)(281),lamdaOut => P(4)(265));
F5266: entity F port map(lamdaA => P(5)(266),lamdaB => P(5)(282),lamdaOut => P(4)(266));
F5267: entity F port map(lamdaA => P(5)(267),lamdaB => P(5)(283),lamdaOut => P(4)(267));
F5268: entity F port map(lamdaA => P(5)(268),lamdaB => P(5)(284),lamdaOut => P(4)(268));
F5269: entity F port map(lamdaA => P(5)(269),lamdaB => P(5)(285),lamdaOut => P(4)(269));
F5270: entity F port map(lamdaA => P(5)(270),lamdaB => P(5)(286),lamdaOut => P(4)(270));
F5271: entity F port map(lamdaA => P(5)(271),lamdaB => P(5)(287),lamdaOut => P(4)(271));
G5272: entity G port map(lamdaA => P(5)(256),lamdaB => P(5)(272),s => s(5)(128),lamdaOut => P(4)(272));
G5273: entity G port map(lamdaA => P(5)(257),lamdaB => P(5)(273),s => s(5)(129),lamdaOut => P(4)(273));
G5274: entity G port map(lamdaA => P(5)(258),lamdaB => P(5)(274),s => s(5)(130),lamdaOut => P(4)(274));
G5275: entity G port map(lamdaA => P(5)(259),lamdaB => P(5)(275),s => s(5)(131),lamdaOut => P(4)(275));
G5276: entity G port map(lamdaA => P(5)(260),lamdaB => P(5)(276),s => s(5)(132),lamdaOut => P(4)(276));
G5277: entity G port map(lamdaA => P(5)(261),lamdaB => P(5)(277),s => s(5)(133),lamdaOut => P(4)(277));
G5278: entity G port map(lamdaA => P(5)(262),lamdaB => P(5)(278),s => s(5)(134),lamdaOut => P(4)(278));
G5279: entity G port map(lamdaA => P(5)(263),lamdaB => P(5)(279),s => s(5)(135),lamdaOut => P(4)(279));
G5280: entity G port map(lamdaA => P(5)(264),lamdaB => P(5)(280),s => s(5)(136),lamdaOut => P(4)(280));
G5281: entity G port map(lamdaA => P(5)(265),lamdaB => P(5)(281),s => s(5)(137),lamdaOut => P(4)(281));
G5282: entity G port map(lamdaA => P(5)(266),lamdaB => P(5)(282),s => s(5)(138),lamdaOut => P(4)(282));
G5283: entity G port map(lamdaA => P(5)(267),lamdaB => P(5)(283),s => s(5)(139),lamdaOut => P(4)(283));
G5284: entity G port map(lamdaA => P(5)(268),lamdaB => P(5)(284),s => s(5)(140),lamdaOut => P(4)(284));
G5285: entity G port map(lamdaA => P(5)(269),lamdaB => P(5)(285),s => s(5)(141),lamdaOut => P(4)(285));
G5286: entity G port map(lamdaA => P(5)(270),lamdaB => P(5)(286),s => s(5)(142),lamdaOut => P(4)(286));
G5287: entity G port map(lamdaA => P(5)(271),lamdaB => P(5)(287),s => s(5)(143),lamdaOut => P(4)(287));
F5288: entity F port map(lamdaA => P(5)(288),lamdaB => P(5)(304),lamdaOut => P(4)(288));
F5289: entity F port map(lamdaA => P(5)(289),lamdaB => P(5)(305),lamdaOut => P(4)(289));
F5290: entity F port map(lamdaA => P(5)(290),lamdaB => P(5)(306),lamdaOut => P(4)(290));
F5291: entity F port map(lamdaA => P(5)(291),lamdaB => P(5)(307),lamdaOut => P(4)(291));
F5292: entity F port map(lamdaA => P(5)(292),lamdaB => P(5)(308),lamdaOut => P(4)(292));
F5293: entity F port map(lamdaA => P(5)(293),lamdaB => P(5)(309),lamdaOut => P(4)(293));
F5294: entity F port map(lamdaA => P(5)(294),lamdaB => P(5)(310),lamdaOut => P(4)(294));
F5295: entity F port map(lamdaA => P(5)(295),lamdaB => P(5)(311),lamdaOut => P(4)(295));
F5296: entity F port map(lamdaA => P(5)(296),lamdaB => P(5)(312),lamdaOut => P(4)(296));
F5297: entity F port map(lamdaA => P(5)(297),lamdaB => P(5)(313),lamdaOut => P(4)(297));
F5298: entity F port map(lamdaA => P(5)(298),lamdaB => P(5)(314),lamdaOut => P(4)(298));
F5299: entity F port map(lamdaA => P(5)(299),lamdaB => P(5)(315),lamdaOut => P(4)(299));
F5300: entity F port map(lamdaA => P(5)(300),lamdaB => P(5)(316),lamdaOut => P(4)(300));
F5301: entity F port map(lamdaA => P(5)(301),lamdaB => P(5)(317),lamdaOut => P(4)(301));
F5302: entity F port map(lamdaA => P(5)(302),lamdaB => P(5)(318),lamdaOut => P(4)(302));
F5303: entity F port map(lamdaA => P(5)(303),lamdaB => P(5)(319),lamdaOut => P(4)(303));
G5304: entity G port map(lamdaA => P(5)(288),lamdaB => P(5)(304),s => s(5)(144),lamdaOut => P(4)(304));
G5305: entity G port map(lamdaA => P(5)(289),lamdaB => P(5)(305),s => s(5)(145),lamdaOut => P(4)(305));
G5306: entity G port map(lamdaA => P(5)(290),lamdaB => P(5)(306),s => s(5)(146),lamdaOut => P(4)(306));
G5307: entity G port map(lamdaA => P(5)(291),lamdaB => P(5)(307),s => s(5)(147),lamdaOut => P(4)(307));
G5308: entity G port map(lamdaA => P(5)(292),lamdaB => P(5)(308),s => s(5)(148),lamdaOut => P(4)(308));
G5309: entity G port map(lamdaA => P(5)(293),lamdaB => P(5)(309),s => s(5)(149),lamdaOut => P(4)(309));
G5310: entity G port map(lamdaA => P(5)(294),lamdaB => P(5)(310),s => s(5)(150),lamdaOut => P(4)(310));
G5311: entity G port map(lamdaA => P(5)(295),lamdaB => P(5)(311),s => s(5)(151),lamdaOut => P(4)(311));
G5312: entity G port map(lamdaA => P(5)(296),lamdaB => P(5)(312),s => s(5)(152),lamdaOut => P(4)(312));
G5313: entity G port map(lamdaA => P(5)(297),lamdaB => P(5)(313),s => s(5)(153),lamdaOut => P(4)(313));
G5314: entity G port map(lamdaA => P(5)(298),lamdaB => P(5)(314),s => s(5)(154),lamdaOut => P(4)(314));
G5315: entity G port map(lamdaA => P(5)(299),lamdaB => P(5)(315),s => s(5)(155),lamdaOut => P(4)(315));
G5316: entity G port map(lamdaA => P(5)(300),lamdaB => P(5)(316),s => s(5)(156),lamdaOut => P(4)(316));
G5317: entity G port map(lamdaA => P(5)(301),lamdaB => P(5)(317),s => s(5)(157),lamdaOut => P(4)(317));
G5318: entity G port map(lamdaA => P(5)(302),lamdaB => P(5)(318),s => s(5)(158),lamdaOut => P(4)(318));
G5319: entity G port map(lamdaA => P(5)(303),lamdaB => P(5)(319),s => s(5)(159),lamdaOut => P(4)(319));
F5320: entity F port map(lamdaA => P(5)(320),lamdaB => P(5)(336),lamdaOut => P(4)(320));
F5321: entity F port map(lamdaA => P(5)(321),lamdaB => P(5)(337),lamdaOut => P(4)(321));
F5322: entity F port map(lamdaA => P(5)(322),lamdaB => P(5)(338),lamdaOut => P(4)(322));
F5323: entity F port map(lamdaA => P(5)(323),lamdaB => P(5)(339),lamdaOut => P(4)(323));
F5324: entity F port map(lamdaA => P(5)(324),lamdaB => P(5)(340),lamdaOut => P(4)(324));
F5325: entity F port map(lamdaA => P(5)(325),lamdaB => P(5)(341),lamdaOut => P(4)(325));
F5326: entity F port map(lamdaA => P(5)(326),lamdaB => P(5)(342),lamdaOut => P(4)(326));
F5327: entity F port map(lamdaA => P(5)(327),lamdaB => P(5)(343),lamdaOut => P(4)(327));
F5328: entity F port map(lamdaA => P(5)(328),lamdaB => P(5)(344),lamdaOut => P(4)(328));
F5329: entity F port map(lamdaA => P(5)(329),lamdaB => P(5)(345),lamdaOut => P(4)(329));
F5330: entity F port map(lamdaA => P(5)(330),lamdaB => P(5)(346),lamdaOut => P(4)(330));
F5331: entity F port map(lamdaA => P(5)(331),lamdaB => P(5)(347),lamdaOut => P(4)(331));
F5332: entity F port map(lamdaA => P(5)(332),lamdaB => P(5)(348),lamdaOut => P(4)(332));
F5333: entity F port map(lamdaA => P(5)(333),lamdaB => P(5)(349),lamdaOut => P(4)(333));
F5334: entity F port map(lamdaA => P(5)(334),lamdaB => P(5)(350),lamdaOut => P(4)(334));
F5335: entity F port map(lamdaA => P(5)(335),lamdaB => P(5)(351),lamdaOut => P(4)(335));
G5336: entity G port map(lamdaA => P(5)(320),lamdaB => P(5)(336),s => s(5)(160),lamdaOut => P(4)(336));
G5337: entity G port map(lamdaA => P(5)(321),lamdaB => P(5)(337),s => s(5)(161),lamdaOut => P(4)(337));
G5338: entity G port map(lamdaA => P(5)(322),lamdaB => P(5)(338),s => s(5)(162),lamdaOut => P(4)(338));
G5339: entity G port map(lamdaA => P(5)(323),lamdaB => P(5)(339),s => s(5)(163),lamdaOut => P(4)(339));
G5340: entity G port map(lamdaA => P(5)(324),lamdaB => P(5)(340),s => s(5)(164),lamdaOut => P(4)(340));
G5341: entity G port map(lamdaA => P(5)(325),lamdaB => P(5)(341),s => s(5)(165),lamdaOut => P(4)(341));
G5342: entity G port map(lamdaA => P(5)(326),lamdaB => P(5)(342),s => s(5)(166),lamdaOut => P(4)(342));
G5343: entity G port map(lamdaA => P(5)(327),lamdaB => P(5)(343),s => s(5)(167),lamdaOut => P(4)(343));
G5344: entity G port map(lamdaA => P(5)(328),lamdaB => P(5)(344),s => s(5)(168),lamdaOut => P(4)(344));
G5345: entity G port map(lamdaA => P(5)(329),lamdaB => P(5)(345),s => s(5)(169),lamdaOut => P(4)(345));
G5346: entity G port map(lamdaA => P(5)(330),lamdaB => P(5)(346),s => s(5)(170),lamdaOut => P(4)(346));
G5347: entity G port map(lamdaA => P(5)(331),lamdaB => P(5)(347),s => s(5)(171),lamdaOut => P(4)(347));
G5348: entity G port map(lamdaA => P(5)(332),lamdaB => P(5)(348),s => s(5)(172),lamdaOut => P(4)(348));
G5349: entity G port map(lamdaA => P(5)(333),lamdaB => P(5)(349),s => s(5)(173),lamdaOut => P(4)(349));
G5350: entity G port map(lamdaA => P(5)(334),lamdaB => P(5)(350),s => s(5)(174),lamdaOut => P(4)(350));
G5351: entity G port map(lamdaA => P(5)(335),lamdaB => P(5)(351),s => s(5)(175),lamdaOut => P(4)(351));
F5352: entity F port map(lamdaA => P(5)(352),lamdaB => P(5)(368),lamdaOut => P(4)(352));
F5353: entity F port map(lamdaA => P(5)(353),lamdaB => P(5)(369),lamdaOut => P(4)(353));
F5354: entity F port map(lamdaA => P(5)(354),lamdaB => P(5)(370),lamdaOut => P(4)(354));
F5355: entity F port map(lamdaA => P(5)(355),lamdaB => P(5)(371),lamdaOut => P(4)(355));
F5356: entity F port map(lamdaA => P(5)(356),lamdaB => P(5)(372),lamdaOut => P(4)(356));
F5357: entity F port map(lamdaA => P(5)(357),lamdaB => P(5)(373),lamdaOut => P(4)(357));
F5358: entity F port map(lamdaA => P(5)(358),lamdaB => P(5)(374),lamdaOut => P(4)(358));
F5359: entity F port map(lamdaA => P(5)(359),lamdaB => P(5)(375),lamdaOut => P(4)(359));
F5360: entity F port map(lamdaA => P(5)(360),lamdaB => P(5)(376),lamdaOut => P(4)(360));
F5361: entity F port map(lamdaA => P(5)(361),lamdaB => P(5)(377),lamdaOut => P(4)(361));
F5362: entity F port map(lamdaA => P(5)(362),lamdaB => P(5)(378),lamdaOut => P(4)(362));
F5363: entity F port map(lamdaA => P(5)(363),lamdaB => P(5)(379),lamdaOut => P(4)(363));
F5364: entity F port map(lamdaA => P(5)(364),lamdaB => P(5)(380),lamdaOut => P(4)(364));
F5365: entity F port map(lamdaA => P(5)(365),lamdaB => P(5)(381),lamdaOut => P(4)(365));
F5366: entity F port map(lamdaA => P(5)(366),lamdaB => P(5)(382),lamdaOut => P(4)(366));
F5367: entity F port map(lamdaA => P(5)(367),lamdaB => P(5)(383),lamdaOut => P(4)(367));
G5368: entity G port map(lamdaA => P(5)(352),lamdaB => P(5)(368),s => s(5)(176),lamdaOut => P(4)(368));
G5369: entity G port map(lamdaA => P(5)(353),lamdaB => P(5)(369),s => s(5)(177),lamdaOut => P(4)(369));
G5370: entity G port map(lamdaA => P(5)(354),lamdaB => P(5)(370),s => s(5)(178),lamdaOut => P(4)(370));
G5371: entity G port map(lamdaA => P(5)(355),lamdaB => P(5)(371),s => s(5)(179),lamdaOut => P(4)(371));
G5372: entity G port map(lamdaA => P(5)(356),lamdaB => P(5)(372),s => s(5)(180),lamdaOut => P(4)(372));
G5373: entity G port map(lamdaA => P(5)(357),lamdaB => P(5)(373),s => s(5)(181),lamdaOut => P(4)(373));
G5374: entity G port map(lamdaA => P(5)(358),lamdaB => P(5)(374),s => s(5)(182),lamdaOut => P(4)(374));
G5375: entity G port map(lamdaA => P(5)(359),lamdaB => P(5)(375),s => s(5)(183),lamdaOut => P(4)(375));
G5376: entity G port map(lamdaA => P(5)(360),lamdaB => P(5)(376),s => s(5)(184),lamdaOut => P(4)(376));
G5377: entity G port map(lamdaA => P(5)(361),lamdaB => P(5)(377),s => s(5)(185),lamdaOut => P(4)(377));
G5378: entity G port map(lamdaA => P(5)(362),lamdaB => P(5)(378),s => s(5)(186),lamdaOut => P(4)(378));
G5379: entity G port map(lamdaA => P(5)(363),lamdaB => P(5)(379),s => s(5)(187),lamdaOut => P(4)(379));
G5380: entity G port map(lamdaA => P(5)(364),lamdaB => P(5)(380),s => s(5)(188),lamdaOut => P(4)(380));
G5381: entity G port map(lamdaA => P(5)(365),lamdaB => P(5)(381),s => s(5)(189),lamdaOut => P(4)(381));
G5382: entity G port map(lamdaA => P(5)(366),lamdaB => P(5)(382),s => s(5)(190),lamdaOut => P(4)(382));
G5383: entity G port map(lamdaA => P(5)(367),lamdaB => P(5)(383),s => s(5)(191),lamdaOut => P(4)(383));
F5384: entity F port map(lamdaA => P(5)(384),lamdaB => P(5)(400),lamdaOut => P(4)(384));
F5385: entity F port map(lamdaA => P(5)(385),lamdaB => P(5)(401),lamdaOut => P(4)(385));
F5386: entity F port map(lamdaA => P(5)(386),lamdaB => P(5)(402),lamdaOut => P(4)(386));
F5387: entity F port map(lamdaA => P(5)(387),lamdaB => P(5)(403),lamdaOut => P(4)(387));
F5388: entity F port map(lamdaA => P(5)(388),lamdaB => P(5)(404),lamdaOut => P(4)(388));
F5389: entity F port map(lamdaA => P(5)(389),lamdaB => P(5)(405),lamdaOut => P(4)(389));
F5390: entity F port map(lamdaA => P(5)(390),lamdaB => P(5)(406),lamdaOut => P(4)(390));
F5391: entity F port map(lamdaA => P(5)(391),lamdaB => P(5)(407),lamdaOut => P(4)(391));
F5392: entity F port map(lamdaA => P(5)(392),lamdaB => P(5)(408),lamdaOut => P(4)(392));
F5393: entity F port map(lamdaA => P(5)(393),lamdaB => P(5)(409),lamdaOut => P(4)(393));
F5394: entity F port map(lamdaA => P(5)(394),lamdaB => P(5)(410),lamdaOut => P(4)(394));
F5395: entity F port map(lamdaA => P(5)(395),lamdaB => P(5)(411),lamdaOut => P(4)(395));
F5396: entity F port map(lamdaA => P(5)(396),lamdaB => P(5)(412),lamdaOut => P(4)(396));
F5397: entity F port map(lamdaA => P(5)(397),lamdaB => P(5)(413),lamdaOut => P(4)(397));
F5398: entity F port map(lamdaA => P(5)(398),lamdaB => P(5)(414),lamdaOut => P(4)(398));
F5399: entity F port map(lamdaA => P(5)(399),lamdaB => P(5)(415),lamdaOut => P(4)(399));
G5400: entity G port map(lamdaA => P(5)(384),lamdaB => P(5)(400),s => s(5)(192),lamdaOut => P(4)(400));
G5401: entity G port map(lamdaA => P(5)(385),lamdaB => P(5)(401),s => s(5)(193),lamdaOut => P(4)(401));
G5402: entity G port map(lamdaA => P(5)(386),lamdaB => P(5)(402),s => s(5)(194),lamdaOut => P(4)(402));
G5403: entity G port map(lamdaA => P(5)(387),lamdaB => P(5)(403),s => s(5)(195),lamdaOut => P(4)(403));
G5404: entity G port map(lamdaA => P(5)(388),lamdaB => P(5)(404),s => s(5)(196),lamdaOut => P(4)(404));
G5405: entity G port map(lamdaA => P(5)(389),lamdaB => P(5)(405),s => s(5)(197),lamdaOut => P(4)(405));
G5406: entity G port map(lamdaA => P(5)(390),lamdaB => P(5)(406),s => s(5)(198),lamdaOut => P(4)(406));
G5407: entity G port map(lamdaA => P(5)(391),lamdaB => P(5)(407),s => s(5)(199),lamdaOut => P(4)(407));
G5408: entity G port map(lamdaA => P(5)(392),lamdaB => P(5)(408),s => s(5)(200),lamdaOut => P(4)(408));
G5409: entity G port map(lamdaA => P(5)(393),lamdaB => P(5)(409),s => s(5)(201),lamdaOut => P(4)(409));
G5410: entity G port map(lamdaA => P(5)(394),lamdaB => P(5)(410),s => s(5)(202),lamdaOut => P(4)(410));
G5411: entity G port map(lamdaA => P(5)(395),lamdaB => P(5)(411),s => s(5)(203),lamdaOut => P(4)(411));
G5412: entity G port map(lamdaA => P(5)(396),lamdaB => P(5)(412),s => s(5)(204),lamdaOut => P(4)(412));
G5413: entity G port map(lamdaA => P(5)(397),lamdaB => P(5)(413),s => s(5)(205),lamdaOut => P(4)(413));
G5414: entity G port map(lamdaA => P(5)(398),lamdaB => P(5)(414),s => s(5)(206),lamdaOut => P(4)(414));
G5415: entity G port map(lamdaA => P(5)(399),lamdaB => P(5)(415),s => s(5)(207),lamdaOut => P(4)(415));
F5416: entity F port map(lamdaA => P(5)(416),lamdaB => P(5)(432),lamdaOut => P(4)(416));
F5417: entity F port map(lamdaA => P(5)(417),lamdaB => P(5)(433),lamdaOut => P(4)(417));
F5418: entity F port map(lamdaA => P(5)(418),lamdaB => P(5)(434),lamdaOut => P(4)(418));
F5419: entity F port map(lamdaA => P(5)(419),lamdaB => P(5)(435),lamdaOut => P(4)(419));
F5420: entity F port map(lamdaA => P(5)(420),lamdaB => P(5)(436),lamdaOut => P(4)(420));
F5421: entity F port map(lamdaA => P(5)(421),lamdaB => P(5)(437),lamdaOut => P(4)(421));
F5422: entity F port map(lamdaA => P(5)(422),lamdaB => P(5)(438),lamdaOut => P(4)(422));
F5423: entity F port map(lamdaA => P(5)(423),lamdaB => P(5)(439),lamdaOut => P(4)(423));
F5424: entity F port map(lamdaA => P(5)(424),lamdaB => P(5)(440),lamdaOut => P(4)(424));
F5425: entity F port map(lamdaA => P(5)(425),lamdaB => P(5)(441),lamdaOut => P(4)(425));
F5426: entity F port map(lamdaA => P(5)(426),lamdaB => P(5)(442),lamdaOut => P(4)(426));
F5427: entity F port map(lamdaA => P(5)(427),lamdaB => P(5)(443),lamdaOut => P(4)(427));
F5428: entity F port map(lamdaA => P(5)(428),lamdaB => P(5)(444),lamdaOut => P(4)(428));
F5429: entity F port map(lamdaA => P(5)(429),lamdaB => P(5)(445),lamdaOut => P(4)(429));
F5430: entity F port map(lamdaA => P(5)(430),lamdaB => P(5)(446),lamdaOut => P(4)(430));
F5431: entity F port map(lamdaA => P(5)(431),lamdaB => P(5)(447),lamdaOut => P(4)(431));
G5432: entity G port map(lamdaA => P(5)(416),lamdaB => P(5)(432),s => s(5)(208),lamdaOut => P(4)(432));
G5433: entity G port map(lamdaA => P(5)(417),lamdaB => P(5)(433),s => s(5)(209),lamdaOut => P(4)(433));
G5434: entity G port map(lamdaA => P(5)(418),lamdaB => P(5)(434),s => s(5)(210),lamdaOut => P(4)(434));
G5435: entity G port map(lamdaA => P(5)(419),lamdaB => P(5)(435),s => s(5)(211),lamdaOut => P(4)(435));
G5436: entity G port map(lamdaA => P(5)(420),lamdaB => P(5)(436),s => s(5)(212),lamdaOut => P(4)(436));
G5437: entity G port map(lamdaA => P(5)(421),lamdaB => P(5)(437),s => s(5)(213),lamdaOut => P(4)(437));
G5438: entity G port map(lamdaA => P(5)(422),lamdaB => P(5)(438),s => s(5)(214),lamdaOut => P(4)(438));
G5439: entity G port map(lamdaA => P(5)(423),lamdaB => P(5)(439),s => s(5)(215),lamdaOut => P(4)(439));
G5440: entity G port map(lamdaA => P(5)(424),lamdaB => P(5)(440),s => s(5)(216),lamdaOut => P(4)(440));
G5441: entity G port map(lamdaA => P(5)(425),lamdaB => P(5)(441),s => s(5)(217),lamdaOut => P(4)(441));
G5442: entity G port map(lamdaA => P(5)(426),lamdaB => P(5)(442),s => s(5)(218),lamdaOut => P(4)(442));
G5443: entity G port map(lamdaA => P(5)(427),lamdaB => P(5)(443),s => s(5)(219),lamdaOut => P(4)(443));
G5444: entity G port map(lamdaA => P(5)(428),lamdaB => P(5)(444),s => s(5)(220),lamdaOut => P(4)(444));
G5445: entity G port map(lamdaA => P(5)(429),lamdaB => P(5)(445),s => s(5)(221),lamdaOut => P(4)(445));
G5446: entity G port map(lamdaA => P(5)(430),lamdaB => P(5)(446),s => s(5)(222),lamdaOut => P(4)(446));
G5447: entity G port map(lamdaA => P(5)(431),lamdaB => P(5)(447),s => s(5)(223),lamdaOut => P(4)(447));
F5448: entity F port map(lamdaA => P(5)(448),lamdaB => P(5)(464),lamdaOut => P(4)(448));
F5449: entity F port map(lamdaA => P(5)(449),lamdaB => P(5)(465),lamdaOut => P(4)(449));
F5450: entity F port map(lamdaA => P(5)(450),lamdaB => P(5)(466),lamdaOut => P(4)(450));
F5451: entity F port map(lamdaA => P(5)(451),lamdaB => P(5)(467),lamdaOut => P(4)(451));
F5452: entity F port map(lamdaA => P(5)(452),lamdaB => P(5)(468),lamdaOut => P(4)(452));
F5453: entity F port map(lamdaA => P(5)(453),lamdaB => P(5)(469),lamdaOut => P(4)(453));
F5454: entity F port map(lamdaA => P(5)(454),lamdaB => P(5)(470),lamdaOut => P(4)(454));
F5455: entity F port map(lamdaA => P(5)(455),lamdaB => P(5)(471),lamdaOut => P(4)(455));
F5456: entity F port map(lamdaA => P(5)(456),lamdaB => P(5)(472),lamdaOut => P(4)(456));
F5457: entity F port map(lamdaA => P(5)(457),lamdaB => P(5)(473),lamdaOut => P(4)(457));
F5458: entity F port map(lamdaA => P(5)(458),lamdaB => P(5)(474),lamdaOut => P(4)(458));
F5459: entity F port map(lamdaA => P(5)(459),lamdaB => P(5)(475),lamdaOut => P(4)(459));
F5460: entity F port map(lamdaA => P(5)(460),lamdaB => P(5)(476),lamdaOut => P(4)(460));
F5461: entity F port map(lamdaA => P(5)(461),lamdaB => P(5)(477),lamdaOut => P(4)(461));
F5462: entity F port map(lamdaA => P(5)(462),lamdaB => P(5)(478),lamdaOut => P(4)(462));
F5463: entity F port map(lamdaA => P(5)(463),lamdaB => P(5)(479),lamdaOut => P(4)(463));
G5464: entity G port map(lamdaA => P(5)(448),lamdaB => P(5)(464),s => s(5)(224),lamdaOut => P(4)(464));
G5465: entity G port map(lamdaA => P(5)(449),lamdaB => P(5)(465),s => s(5)(225),lamdaOut => P(4)(465));
G5466: entity G port map(lamdaA => P(5)(450),lamdaB => P(5)(466),s => s(5)(226),lamdaOut => P(4)(466));
G5467: entity G port map(lamdaA => P(5)(451),lamdaB => P(5)(467),s => s(5)(227),lamdaOut => P(4)(467));
G5468: entity G port map(lamdaA => P(5)(452),lamdaB => P(5)(468),s => s(5)(228),lamdaOut => P(4)(468));
G5469: entity G port map(lamdaA => P(5)(453),lamdaB => P(5)(469),s => s(5)(229),lamdaOut => P(4)(469));
G5470: entity G port map(lamdaA => P(5)(454),lamdaB => P(5)(470),s => s(5)(230),lamdaOut => P(4)(470));
G5471: entity G port map(lamdaA => P(5)(455),lamdaB => P(5)(471),s => s(5)(231),lamdaOut => P(4)(471));
G5472: entity G port map(lamdaA => P(5)(456),lamdaB => P(5)(472),s => s(5)(232),lamdaOut => P(4)(472));
G5473: entity G port map(lamdaA => P(5)(457),lamdaB => P(5)(473),s => s(5)(233),lamdaOut => P(4)(473));
G5474: entity G port map(lamdaA => P(5)(458),lamdaB => P(5)(474),s => s(5)(234),lamdaOut => P(4)(474));
G5475: entity G port map(lamdaA => P(5)(459),lamdaB => P(5)(475),s => s(5)(235),lamdaOut => P(4)(475));
G5476: entity G port map(lamdaA => P(5)(460),lamdaB => P(5)(476),s => s(5)(236),lamdaOut => P(4)(476));
G5477: entity G port map(lamdaA => P(5)(461),lamdaB => P(5)(477),s => s(5)(237),lamdaOut => P(4)(477));
G5478: entity G port map(lamdaA => P(5)(462),lamdaB => P(5)(478),s => s(5)(238),lamdaOut => P(4)(478));
G5479: entity G port map(lamdaA => P(5)(463),lamdaB => P(5)(479),s => s(5)(239),lamdaOut => P(4)(479));
F5480: entity F port map(lamdaA => P(5)(480),lamdaB => P(5)(496),lamdaOut => P(4)(480));
F5481: entity F port map(lamdaA => P(5)(481),lamdaB => P(5)(497),lamdaOut => P(4)(481));
F5482: entity F port map(lamdaA => P(5)(482),lamdaB => P(5)(498),lamdaOut => P(4)(482));
F5483: entity F port map(lamdaA => P(5)(483),lamdaB => P(5)(499),lamdaOut => P(4)(483));
F5484: entity F port map(lamdaA => P(5)(484),lamdaB => P(5)(500),lamdaOut => P(4)(484));
F5485: entity F port map(lamdaA => P(5)(485),lamdaB => P(5)(501),lamdaOut => P(4)(485));
F5486: entity F port map(lamdaA => P(5)(486),lamdaB => P(5)(502),lamdaOut => P(4)(486));
F5487: entity F port map(lamdaA => P(5)(487),lamdaB => P(5)(503),lamdaOut => P(4)(487));
F5488: entity F port map(lamdaA => P(5)(488),lamdaB => P(5)(504),lamdaOut => P(4)(488));
F5489: entity F port map(lamdaA => P(5)(489),lamdaB => P(5)(505),lamdaOut => P(4)(489));
F5490: entity F port map(lamdaA => P(5)(490),lamdaB => P(5)(506),lamdaOut => P(4)(490));
F5491: entity F port map(lamdaA => P(5)(491),lamdaB => P(5)(507),lamdaOut => P(4)(491));
F5492: entity F port map(lamdaA => P(5)(492),lamdaB => P(5)(508),lamdaOut => P(4)(492));
F5493: entity F port map(lamdaA => P(5)(493),lamdaB => P(5)(509),lamdaOut => P(4)(493));
F5494: entity F port map(lamdaA => P(5)(494),lamdaB => P(5)(510),lamdaOut => P(4)(494));
F5495: entity F port map(lamdaA => P(5)(495),lamdaB => P(5)(511),lamdaOut => P(4)(495));
G5496: entity G port map(lamdaA => P(5)(480),lamdaB => P(5)(496),s => s(5)(240),lamdaOut => P(4)(496));
G5497: entity G port map(lamdaA => P(5)(481),lamdaB => P(5)(497),s => s(5)(241),lamdaOut => P(4)(497));
G5498: entity G port map(lamdaA => P(5)(482),lamdaB => P(5)(498),s => s(5)(242),lamdaOut => P(4)(498));
G5499: entity G port map(lamdaA => P(5)(483),lamdaB => P(5)(499),s => s(5)(243),lamdaOut => P(4)(499));
G5500: entity G port map(lamdaA => P(5)(484),lamdaB => P(5)(500),s => s(5)(244),lamdaOut => P(4)(500));
G5501: entity G port map(lamdaA => P(5)(485),lamdaB => P(5)(501),s => s(5)(245),lamdaOut => P(4)(501));
G5502: entity G port map(lamdaA => P(5)(486),lamdaB => P(5)(502),s => s(5)(246),lamdaOut => P(4)(502));
G5503: entity G port map(lamdaA => P(5)(487),lamdaB => P(5)(503),s => s(5)(247),lamdaOut => P(4)(503));
G5504: entity G port map(lamdaA => P(5)(488),lamdaB => P(5)(504),s => s(5)(248),lamdaOut => P(4)(504));
G5505: entity G port map(lamdaA => P(5)(489),lamdaB => P(5)(505),s => s(5)(249),lamdaOut => P(4)(505));
G5506: entity G port map(lamdaA => P(5)(490),lamdaB => P(5)(506),s => s(5)(250),lamdaOut => P(4)(506));
G5507: entity G port map(lamdaA => P(5)(491),lamdaB => P(5)(507),s => s(5)(251),lamdaOut => P(4)(507));
G5508: entity G port map(lamdaA => P(5)(492),lamdaB => P(5)(508),s => s(5)(252),lamdaOut => P(4)(508));
G5509: entity G port map(lamdaA => P(5)(493),lamdaB => P(5)(509),s => s(5)(253),lamdaOut => P(4)(509));
G5510: entity G port map(lamdaA => P(5)(494),lamdaB => P(5)(510),s => s(5)(254),lamdaOut => P(4)(510));
G5511: entity G port map(lamdaA => P(5)(495),lamdaB => P(5)(511),s => s(5)(255),lamdaOut => P(4)(511));
-- STAGE 4
F40: entity F port map(lamdaA => P(4)(0),lamdaB => P(4)(32),lamdaOut => P(3)(0));
F41: entity F port map(lamdaA => P(4)(1),lamdaB => P(4)(33),lamdaOut => P(3)(1));
F42: entity F port map(lamdaA => P(4)(2),lamdaB => P(4)(34),lamdaOut => P(3)(2));
F43: entity F port map(lamdaA => P(4)(3),lamdaB => P(4)(35),lamdaOut => P(3)(3));
F44: entity F port map(lamdaA => P(4)(4),lamdaB => P(4)(36),lamdaOut => P(3)(4));
F45: entity F port map(lamdaA => P(4)(5),lamdaB => P(4)(37),lamdaOut => P(3)(5));
F46: entity F port map(lamdaA => P(4)(6),lamdaB => P(4)(38),lamdaOut => P(3)(6));
F47: entity F port map(lamdaA => P(4)(7),lamdaB => P(4)(39),lamdaOut => P(3)(7));
F48: entity F port map(lamdaA => P(4)(8),lamdaB => P(4)(40),lamdaOut => P(3)(8));
F49: entity F port map(lamdaA => P(4)(9),lamdaB => P(4)(41),lamdaOut => P(3)(9));
F410: entity F port map(lamdaA => P(4)(10),lamdaB => P(4)(42),lamdaOut => P(3)(10));
F411: entity F port map(lamdaA => P(4)(11),lamdaB => P(4)(43),lamdaOut => P(3)(11));
F412: entity F port map(lamdaA => P(4)(12),lamdaB => P(4)(44),lamdaOut => P(3)(12));
F413: entity F port map(lamdaA => P(4)(13),lamdaB => P(4)(45),lamdaOut => P(3)(13));
F414: entity F port map(lamdaA => P(4)(14),lamdaB => P(4)(46),lamdaOut => P(3)(14));
F415: entity F port map(lamdaA => P(4)(15),lamdaB => P(4)(47),lamdaOut => P(3)(15));
F416: entity F port map(lamdaA => P(4)(16),lamdaB => P(4)(48),lamdaOut => P(3)(16));
F417: entity F port map(lamdaA => P(4)(17),lamdaB => P(4)(49),lamdaOut => P(3)(17));
F418: entity F port map(lamdaA => P(4)(18),lamdaB => P(4)(50),lamdaOut => P(3)(18));
F419: entity F port map(lamdaA => P(4)(19),lamdaB => P(4)(51),lamdaOut => P(3)(19));
F420: entity F port map(lamdaA => P(4)(20),lamdaB => P(4)(52),lamdaOut => P(3)(20));
F421: entity F port map(lamdaA => P(4)(21),lamdaB => P(4)(53),lamdaOut => P(3)(21));
F422: entity F port map(lamdaA => P(4)(22),lamdaB => P(4)(54),lamdaOut => P(3)(22));
F423: entity F port map(lamdaA => P(4)(23),lamdaB => P(4)(55),lamdaOut => P(3)(23));
F424: entity F port map(lamdaA => P(4)(24),lamdaB => P(4)(56),lamdaOut => P(3)(24));
F425: entity F port map(lamdaA => P(4)(25),lamdaB => P(4)(57),lamdaOut => P(3)(25));
F426: entity F port map(lamdaA => P(4)(26),lamdaB => P(4)(58),lamdaOut => P(3)(26));
F427: entity F port map(lamdaA => P(4)(27),lamdaB => P(4)(59),lamdaOut => P(3)(27));
F428: entity F port map(lamdaA => P(4)(28),lamdaB => P(4)(60),lamdaOut => P(3)(28));
F429: entity F port map(lamdaA => P(4)(29),lamdaB => P(4)(61),lamdaOut => P(3)(29));
F430: entity F port map(lamdaA => P(4)(30),lamdaB => P(4)(62),lamdaOut => P(3)(30));
F431: entity F port map(lamdaA => P(4)(31),lamdaB => P(4)(63),lamdaOut => P(3)(31));
G432: entity G port map(lamdaA => P(4)(0),lamdaB => P(4)(32),s => s(4)(0),lamdaOut => P(3)(32));
G433: entity G port map(lamdaA => P(4)(1),lamdaB => P(4)(33),s => s(4)(1),lamdaOut => P(3)(33));
G434: entity G port map(lamdaA => P(4)(2),lamdaB => P(4)(34),s => s(4)(2),lamdaOut => P(3)(34));
G435: entity G port map(lamdaA => P(4)(3),lamdaB => P(4)(35),s => s(4)(3),lamdaOut => P(3)(35));
G436: entity G port map(lamdaA => P(4)(4),lamdaB => P(4)(36),s => s(4)(4),lamdaOut => P(3)(36));
G437: entity G port map(lamdaA => P(4)(5),lamdaB => P(4)(37),s => s(4)(5),lamdaOut => P(3)(37));
G438: entity G port map(lamdaA => P(4)(6),lamdaB => P(4)(38),s => s(4)(6),lamdaOut => P(3)(38));
G439: entity G port map(lamdaA => P(4)(7),lamdaB => P(4)(39),s => s(4)(7),lamdaOut => P(3)(39));
G440: entity G port map(lamdaA => P(4)(8),lamdaB => P(4)(40),s => s(4)(8),lamdaOut => P(3)(40));
G441: entity G port map(lamdaA => P(4)(9),lamdaB => P(4)(41),s => s(4)(9),lamdaOut => P(3)(41));
G442: entity G port map(lamdaA => P(4)(10),lamdaB => P(4)(42),s => s(4)(10),lamdaOut => P(3)(42));
G443: entity G port map(lamdaA => P(4)(11),lamdaB => P(4)(43),s => s(4)(11),lamdaOut => P(3)(43));
G444: entity G port map(lamdaA => P(4)(12),lamdaB => P(4)(44),s => s(4)(12),lamdaOut => P(3)(44));
G445: entity G port map(lamdaA => P(4)(13),lamdaB => P(4)(45),s => s(4)(13),lamdaOut => P(3)(45));
G446: entity G port map(lamdaA => P(4)(14),lamdaB => P(4)(46),s => s(4)(14),lamdaOut => P(3)(46));
G447: entity G port map(lamdaA => P(4)(15),lamdaB => P(4)(47),s => s(4)(15),lamdaOut => P(3)(47));
G448: entity G port map(lamdaA => P(4)(16),lamdaB => P(4)(48),s => s(4)(16),lamdaOut => P(3)(48));
G449: entity G port map(lamdaA => P(4)(17),lamdaB => P(4)(49),s => s(4)(17),lamdaOut => P(3)(49));
G450: entity G port map(lamdaA => P(4)(18),lamdaB => P(4)(50),s => s(4)(18),lamdaOut => P(3)(50));
G451: entity G port map(lamdaA => P(4)(19),lamdaB => P(4)(51),s => s(4)(19),lamdaOut => P(3)(51));
G452: entity G port map(lamdaA => P(4)(20),lamdaB => P(4)(52),s => s(4)(20),lamdaOut => P(3)(52));
G453: entity G port map(lamdaA => P(4)(21),lamdaB => P(4)(53),s => s(4)(21),lamdaOut => P(3)(53));
G454: entity G port map(lamdaA => P(4)(22),lamdaB => P(4)(54),s => s(4)(22),lamdaOut => P(3)(54));
G455: entity G port map(lamdaA => P(4)(23),lamdaB => P(4)(55),s => s(4)(23),lamdaOut => P(3)(55));
G456: entity G port map(lamdaA => P(4)(24),lamdaB => P(4)(56),s => s(4)(24),lamdaOut => P(3)(56));
G457: entity G port map(lamdaA => P(4)(25),lamdaB => P(4)(57),s => s(4)(25),lamdaOut => P(3)(57));
G458: entity G port map(lamdaA => P(4)(26),lamdaB => P(4)(58),s => s(4)(26),lamdaOut => P(3)(58));
G459: entity G port map(lamdaA => P(4)(27),lamdaB => P(4)(59),s => s(4)(27),lamdaOut => P(3)(59));
G460: entity G port map(lamdaA => P(4)(28),lamdaB => P(4)(60),s => s(4)(28),lamdaOut => P(3)(60));
G461: entity G port map(lamdaA => P(4)(29),lamdaB => P(4)(61),s => s(4)(29),lamdaOut => P(3)(61));
G462: entity G port map(lamdaA => P(4)(30),lamdaB => P(4)(62),s => s(4)(30),lamdaOut => P(3)(62));
G463: entity G port map(lamdaA => P(4)(31),lamdaB => P(4)(63),s => s(4)(31),lamdaOut => P(3)(63));
F464: entity F port map(lamdaA => P(4)(64),lamdaB => P(4)(96),lamdaOut => P(3)(64));
F465: entity F port map(lamdaA => P(4)(65),lamdaB => P(4)(97),lamdaOut => P(3)(65));
F466: entity F port map(lamdaA => P(4)(66),lamdaB => P(4)(98),lamdaOut => P(3)(66));
F467: entity F port map(lamdaA => P(4)(67),lamdaB => P(4)(99),lamdaOut => P(3)(67));
F468: entity F port map(lamdaA => P(4)(68),lamdaB => P(4)(100),lamdaOut => P(3)(68));
F469: entity F port map(lamdaA => P(4)(69),lamdaB => P(4)(101),lamdaOut => P(3)(69));
F470: entity F port map(lamdaA => P(4)(70),lamdaB => P(4)(102),lamdaOut => P(3)(70));
F471: entity F port map(lamdaA => P(4)(71),lamdaB => P(4)(103),lamdaOut => P(3)(71));
F472: entity F port map(lamdaA => P(4)(72),lamdaB => P(4)(104),lamdaOut => P(3)(72));
F473: entity F port map(lamdaA => P(4)(73),lamdaB => P(4)(105),lamdaOut => P(3)(73));
F474: entity F port map(lamdaA => P(4)(74),lamdaB => P(4)(106),lamdaOut => P(3)(74));
F475: entity F port map(lamdaA => P(4)(75),lamdaB => P(4)(107),lamdaOut => P(3)(75));
F476: entity F port map(lamdaA => P(4)(76),lamdaB => P(4)(108),lamdaOut => P(3)(76));
F477: entity F port map(lamdaA => P(4)(77),lamdaB => P(4)(109),lamdaOut => P(3)(77));
F478: entity F port map(lamdaA => P(4)(78),lamdaB => P(4)(110),lamdaOut => P(3)(78));
F479: entity F port map(lamdaA => P(4)(79),lamdaB => P(4)(111),lamdaOut => P(3)(79));
F480: entity F port map(lamdaA => P(4)(80),lamdaB => P(4)(112),lamdaOut => P(3)(80));
F481: entity F port map(lamdaA => P(4)(81),lamdaB => P(4)(113),lamdaOut => P(3)(81));
F482: entity F port map(lamdaA => P(4)(82),lamdaB => P(4)(114),lamdaOut => P(3)(82));
F483: entity F port map(lamdaA => P(4)(83),lamdaB => P(4)(115),lamdaOut => P(3)(83));
F484: entity F port map(lamdaA => P(4)(84),lamdaB => P(4)(116),lamdaOut => P(3)(84));
F485: entity F port map(lamdaA => P(4)(85),lamdaB => P(4)(117),lamdaOut => P(3)(85));
F486: entity F port map(lamdaA => P(4)(86),lamdaB => P(4)(118),lamdaOut => P(3)(86));
F487: entity F port map(lamdaA => P(4)(87),lamdaB => P(4)(119),lamdaOut => P(3)(87));
F488: entity F port map(lamdaA => P(4)(88),lamdaB => P(4)(120),lamdaOut => P(3)(88));
F489: entity F port map(lamdaA => P(4)(89),lamdaB => P(4)(121),lamdaOut => P(3)(89));
F490: entity F port map(lamdaA => P(4)(90),lamdaB => P(4)(122),lamdaOut => P(3)(90));
F491: entity F port map(lamdaA => P(4)(91),lamdaB => P(4)(123),lamdaOut => P(3)(91));
F492: entity F port map(lamdaA => P(4)(92),lamdaB => P(4)(124),lamdaOut => P(3)(92));
F493: entity F port map(lamdaA => P(4)(93),lamdaB => P(4)(125),lamdaOut => P(3)(93));
F494: entity F port map(lamdaA => P(4)(94),lamdaB => P(4)(126),lamdaOut => P(3)(94));
F495: entity F port map(lamdaA => P(4)(95),lamdaB => P(4)(127),lamdaOut => P(3)(95));
G496: entity G port map(lamdaA => P(4)(64),lamdaB => P(4)(96),s => s(4)(32),lamdaOut => P(3)(96));
G497: entity G port map(lamdaA => P(4)(65),lamdaB => P(4)(97),s => s(4)(33),lamdaOut => P(3)(97));
G498: entity G port map(lamdaA => P(4)(66),lamdaB => P(4)(98),s => s(4)(34),lamdaOut => P(3)(98));
G499: entity G port map(lamdaA => P(4)(67),lamdaB => P(4)(99),s => s(4)(35),lamdaOut => P(3)(99));
G4100: entity G port map(lamdaA => P(4)(68),lamdaB => P(4)(100),s => s(4)(36),lamdaOut => P(3)(100));
G4101: entity G port map(lamdaA => P(4)(69),lamdaB => P(4)(101),s => s(4)(37),lamdaOut => P(3)(101));
G4102: entity G port map(lamdaA => P(4)(70),lamdaB => P(4)(102),s => s(4)(38),lamdaOut => P(3)(102));
G4103: entity G port map(lamdaA => P(4)(71),lamdaB => P(4)(103),s => s(4)(39),lamdaOut => P(3)(103));
G4104: entity G port map(lamdaA => P(4)(72),lamdaB => P(4)(104),s => s(4)(40),lamdaOut => P(3)(104));
G4105: entity G port map(lamdaA => P(4)(73),lamdaB => P(4)(105),s => s(4)(41),lamdaOut => P(3)(105));
G4106: entity G port map(lamdaA => P(4)(74),lamdaB => P(4)(106),s => s(4)(42),lamdaOut => P(3)(106));
G4107: entity G port map(lamdaA => P(4)(75),lamdaB => P(4)(107),s => s(4)(43),lamdaOut => P(3)(107));
G4108: entity G port map(lamdaA => P(4)(76),lamdaB => P(4)(108),s => s(4)(44),lamdaOut => P(3)(108));
G4109: entity G port map(lamdaA => P(4)(77),lamdaB => P(4)(109),s => s(4)(45),lamdaOut => P(3)(109));
G4110: entity G port map(lamdaA => P(4)(78),lamdaB => P(4)(110),s => s(4)(46),lamdaOut => P(3)(110));
G4111: entity G port map(lamdaA => P(4)(79),lamdaB => P(4)(111),s => s(4)(47),lamdaOut => P(3)(111));
G4112: entity G port map(lamdaA => P(4)(80),lamdaB => P(4)(112),s => s(4)(48),lamdaOut => P(3)(112));
G4113: entity G port map(lamdaA => P(4)(81),lamdaB => P(4)(113),s => s(4)(49),lamdaOut => P(3)(113));
G4114: entity G port map(lamdaA => P(4)(82),lamdaB => P(4)(114),s => s(4)(50),lamdaOut => P(3)(114));
G4115: entity G port map(lamdaA => P(4)(83),lamdaB => P(4)(115),s => s(4)(51),lamdaOut => P(3)(115));
G4116: entity G port map(lamdaA => P(4)(84),lamdaB => P(4)(116),s => s(4)(52),lamdaOut => P(3)(116));
G4117: entity G port map(lamdaA => P(4)(85),lamdaB => P(4)(117),s => s(4)(53),lamdaOut => P(3)(117));
G4118: entity G port map(lamdaA => P(4)(86),lamdaB => P(4)(118),s => s(4)(54),lamdaOut => P(3)(118));
G4119: entity G port map(lamdaA => P(4)(87),lamdaB => P(4)(119),s => s(4)(55),lamdaOut => P(3)(119));
G4120: entity G port map(lamdaA => P(4)(88),lamdaB => P(4)(120),s => s(4)(56),lamdaOut => P(3)(120));
G4121: entity G port map(lamdaA => P(4)(89),lamdaB => P(4)(121),s => s(4)(57),lamdaOut => P(3)(121));
G4122: entity G port map(lamdaA => P(4)(90),lamdaB => P(4)(122),s => s(4)(58),lamdaOut => P(3)(122));
G4123: entity G port map(lamdaA => P(4)(91),lamdaB => P(4)(123),s => s(4)(59),lamdaOut => P(3)(123));
G4124: entity G port map(lamdaA => P(4)(92),lamdaB => P(4)(124),s => s(4)(60),lamdaOut => P(3)(124));
G4125: entity G port map(lamdaA => P(4)(93),lamdaB => P(4)(125),s => s(4)(61),lamdaOut => P(3)(125));
G4126: entity G port map(lamdaA => P(4)(94),lamdaB => P(4)(126),s => s(4)(62),lamdaOut => P(3)(126));
G4127: entity G port map(lamdaA => P(4)(95),lamdaB => P(4)(127),s => s(4)(63),lamdaOut => P(3)(127));
F4128: entity F port map(lamdaA => P(4)(128),lamdaB => P(4)(160),lamdaOut => P(3)(128));
F4129: entity F port map(lamdaA => P(4)(129),lamdaB => P(4)(161),lamdaOut => P(3)(129));
F4130: entity F port map(lamdaA => P(4)(130),lamdaB => P(4)(162),lamdaOut => P(3)(130));
F4131: entity F port map(lamdaA => P(4)(131),lamdaB => P(4)(163),lamdaOut => P(3)(131));
F4132: entity F port map(lamdaA => P(4)(132),lamdaB => P(4)(164),lamdaOut => P(3)(132));
F4133: entity F port map(lamdaA => P(4)(133),lamdaB => P(4)(165),lamdaOut => P(3)(133));
F4134: entity F port map(lamdaA => P(4)(134),lamdaB => P(4)(166),lamdaOut => P(3)(134));
F4135: entity F port map(lamdaA => P(4)(135),lamdaB => P(4)(167),lamdaOut => P(3)(135));
F4136: entity F port map(lamdaA => P(4)(136),lamdaB => P(4)(168),lamdaOut => P(3)(136));
F4137: entity F port map(lamdaA => P(4)(137),lamdaB => P(4)(169),lamdaOut => P(3)(137));
F4138: entity F port map(lamdaA => P(4)(138),lamdaB => P(4)(170),lamdaOut => P(3)(138));
F4139: entity F port map(lamdaA => P(4)(139),lamdaB => P(4)(171),lamdaOut => P(3)(139));
F4140: entity F port map(lamdaA => P(4)(140),lamdaB => P(4)(172),lamdaOut => P(3)(140));
F4141: entity F port map(lamdaA => P(4)(141),lamdaB => P(4)(173),lamdaOut => P(3)(141));
F4142: entity F port map(lamdaA => P(4)(142),lamdaB => P(4)(174),lamdaOut => P(3)(142));
F4143: entity F port map(lamdaA => P(4)(143),lamdaB => P(4)(175),lamdaOut => P(3)(143));
F4144: entity F port map(lamdaA => P(4)(144),lamdaB => P(4)(176),lamdaOut => P(3)(144));
F4145: entity F port map(lamdaA => P(4)(145),lamdaB => P(4)(177),lamdaOut => P(3)(145));
F4146: entity F port map(lamdaA => P(4)(146),lamdaB => P(4)(178),lamdaOut => P(3)(146));
F4147: entity F port map(lamdaA => P(4)(147),lamdaB => P(4)(179),lamdaOut => P(3)(147));
F4148: entity F port map(lamdaA => P(4)(148),lamdaB => P(4)(180),lamdaOut => P(3)(148));
F4149: entity F port map(lamdaA => P(4)(149),lamdaB => P(4)(181),lamdaOut => P(3)(149));
F4150: entity F port map(lamdaA => P(4)(150),lamdaB => P(4)(182),lamdaOut => P(3)(150));
F4151: entity F port map(lamdaA => P(4)(151),lamdaB => P(4)(183),lamdaOut => P(3)(151));
F4152: entity F port map(lamdaA => P(4)(152),lamdaB => P(4)(184),lamdaOut => P(3)(152));
F4153: entity F port map(lamdaA => P(4)(153),lamdaB => P(4)(185),lamdaOut => P(3)(153));
F4154: entity F port map(lamdaA => P(4)(154),lamdaB => P(4)(186),lamdaOut => P(3)(154));
F4155: entity F port map(lamdaA => P(4)(155),lamdaB => P(4)(187),lamdaOut => P(3)(155));
F4156: entity F port map(lamdaA => P(4)(156),lamdaB => P(4)(188),lamdaOut => P(3)(156));
F4157: entity F port map(lamdaA => P(4)(157),lamdaB => P(4)(189),lamdaOut => P(3)(157));
F4158: entity F port map(lamdaA => P(4)(158),lamdaB => P(4)(190),lamdaOut => P(3)(158));
F4159: entity F port map(lamdaA => P(4)(159),lamdaB => P(4)(191),lamdaOut => P(3)(159));
G4160: entity G port map(lamdaA => P(4)(128),lamdaB => P(4)(160),s => s(4)(64),lamdaOut => P(3)(160));
G4161: entity G port map(lamdaA => P(4)(129),lamdaB => P(4)(161),s => s(4)(65),lamdaOut => P(3)(161));
G4162: entity G port map(lamdaA => P(4)(130),lamdaB => P(4)(162),s => s(4)(66),lamdaOut => P(3)(162));
G4163: entity G port map(lamdaA => P(4)(131),lamdaB => P(4)(163),s => s(4)(67),lamdaOut => P(3)(163));
G4164: entity G port map(lamdaA => P(4)(132),lamdaB => P(4)(164),s => s(4)(68),lamdaOut => P(3)(164));
G4165: entity G port map(lamdaA => P(4)(133),lamdaB => P(4)(165),s => s(4)(69),lamdaOut => P(3)(165));
G4166: entity G port map(lamdaA => P(4)(134),lamdaB => P(4)(166),s => s(4)(70),lamdaOut => P(3)(166));
G4167: entity G port map(lamdaA => P(4)(135),lamdaB => P(4)(167),s => s(4)(71),lamdaOut => P(3)(167));
G4168: entity G port map(lamdaA => P(4)(136),lamdaB => P(4)(168),s => s(4)(72),lamdaOut => P(3)(168));
G4169: entity G port map(lamdaA => P(4)(137),lamdaB => P(4)(169),s => s(4)(73),lamdaOut => P(3)(169));
G4170: entity G port map(lamdaA => P(4)(138),lamdaB => P(4)(170),s => s(4)(74),lamdaOut => P(3)(170));
G4171: entity G port map(lamdaA => P(4)(139),lamdaB => P(4)(171),s => s(4)(75),lamdaOut => P(3)(171));
G4172: entity G port map(lamdaA => P(4)(140),lamdaB => P(4)(172),s => s(4)(76),lamdaOut => P(3)(172));
G4173: entity G port map(lamdaA => P(4)(141),lamdaB => P(4)(173),s => s(4)(77),lamdaOut => P(3)(173));
G4174: entity G port map(lamdaA => P(4)(142),lamdaB => P(4)(174),s => s(4)(78),lamdaOut => P(3)(174));
G4175: entity G port map(lamdaA => P(4)(143),lamdaB => P(4)(175),s => s(4)(79),lamdaOut => P(3)(175));
G4176: entity G port map(lamdaA => P(4)(144),lamdaB => P(4)(176),s => s(4)(80),lamdaOut => P(3)(176));
G4177: entity G port map(lamdaA => P(4)(145),lamdaB => P(4)(177),s => s(4)(81),lamdaOut => P(3)(177));
G4178: entity G port map(lamdaA => P(4)(146),lamdaB => P(4)(178),s => s(4)(82),lamdaOut => P(3)(178));
G4179: entity G port map(lamdaA => P(4)(147),lamdaB => P(4)(179),s => s(4)(83),lamdaOut => P(3)(179));
G4180: entity G port map(lamdaA => P(4)(148),lamdaB => P(4)(180),s => s(4)(84),lamdaOut => P(3)(180));
G4181: entity G port map(lamdaA => P(4)(149),lamdaB => P(4)(181),s => s(4)(85),lamdaOut => P(3)(181));
G4182: entity G port map(lamdaA => P(4)(150),lamdaB => P(4)(182),s => s(4)(86),lamdaOut => P(3)(182));
G4183: entity G port map(lamdaA => P(4)(151),lamdaB => P(4)(183),s => s(4)(87),lamdaOut => P(3)(183));
G4184: entity G port map(lamdaA => P(4)(152),lamdaB => P(4)(184),s => s(4)(88),lamdaOut => P(3)(184));
G4185: entity G port map(lamdaA => P(4)(153),lamdaB => P(4)(185),s => s(4)(89),lamdaOut => P(3)(185));
G4186: entity G port map(lamdaA => P(4)(154),lamdaB => P(4)(186),s => s(4)(90),lamdaOut => P(3)(186));
G4187: entity G port map(lamdaA => P(4)(155),lamdaB => P(4)(187),s => s(4)(91),lamdaOut => P(3)(187));
G4188: entity G port map(lamdaA => P(4)(156),lamdaB => P(4)(188),s => s(4)(92),lamdaOut => P(3)(188));
G4189: entity G port map(lamdaA => P(4)(157),lamdaB => P(4)(189),s => s(4)(93),lamdaOut => P(3)(189));
G4190: entity G port map(lamdaA => P(4)(158),lamdaB => P(4)(190),s => s(4)(94),lamdaOut => P(3)(190));
G4191: entity G port map(lamdaA => P(4)(159),lamdaB => P(4)(191),s => s(4)(95),lamdaOut => P(3)(191));
F4192: entity F port map(lamdaA => P(4)(192),lamdaB => P(4)(224),lamdaOut => P(3)(192));
F4193: entity F port map(lamdaA => P(4)(193),lamdaB => P(4)(225),lamdaOut => P(3)(193));
F4194: entity F port map(lamdaA => P(4)(194),lamdaB => P(4)(226),lamdaOut => P(3)(194));
F4195: entity F port map(lamdaA => P(4)(195),lamdaB => P(4)(227),lamdaOut => P(3)(195));
F4196: entity F port map(lamdaA => P(4)(196),lamdaB => P(4)(228),lamdaOut => P(3)(196));
F4197: entity F port map(lamdaA => P(4)(197),lamdaB => P(4)(229),lamdaOut => P(3)(197));
F4198: entity F port map(lamdaA => P(4)(198),lamdaB => P(4)(230),lamdaOut => P(3)(198));
F4199: entity F port map(lamdaA => P(4)(199),lamdaB => P(4)(231),lamdaOut => P(3)(199));
F4200: entity F port map(lamdaA => P(4)(200),lamdaB => P(4)(232),lamdaOut => P(3)(200));
F4201: entity F port map(lamdaA => P(4)(201),lamdaB => P(4)(233),lamdaOut => P(3)(201));
F4202: entity F port map(lamdaA => P(4)(202),lamdaB => P(4)(234),lamdaOut => P(3)(202));
F4203: entity F port map(lamdaA => P(4)(203),lamdaB => P(4)(235),lamdaOut => P(3)(203));
F4204: entity F port map(lamdaA => P(4)(204),lamdaB => P(4)(236),lamdaOut => P(3)(204));
F4205: entity F port map(lamdaA => P(4)(205),lamdaB => P(4)(237),lamdaOut => P(3)(205));
F4206: entity F port map(lamdaA => P(4)(206),lamdaB => P(4)(238),lamdaOut => P(3)(206));
F4207: entity F port map(lamdaA => P(4)(207),lamdaB => P(4)(239),lamdaOut => P(3)(207));
F4208: entity F port map(lamdaA => P(4)(208),lamdaB => P(4)(240),lamdaOut => P(3)(208));
F4209: entity F port map(lamdaA => P(4)(209),lamdaB => P(4)(241),lamdaOut => P(3)(209));
F4210: entity F port map(lamdaA => P(4)(210),lamdaB => P(4)(242),lamdaOut => P(3)(210));
F4211: entity F port map(lamdaA => P(4)(211),lamdaB => P(4)(243),lamdaOut => P(3)(211));
F4212: entity F port map(lamdaA => P(4)(212),lamdaB => P(4)(244),lamdaOut => P(3)(212));
F4213: entity F port map(lamdaA => P(4)(213),lamdaB => P(4)(245),lamdaOut => P(3)(213));
F4214: entity F port map(lamdaA => P(4)(214),lamdaB => P(4)(246),lamdaOut => P(3)(214));
F4215: entity F port map(lamdaA => P(4)(215),lamdaB => P(4)(247),lamdaOut => P(3)(215));
F4216: entity F port map(lamdaA => P(4)(216),lamdaB => P(4)(248),lamdaOut => P(3)(216));
F4217: entity F port map(lamdaA => P(4)(217),lamdaB => P(4)(249),lamdaOut => P(3)(217));
F4218: entity F port map(lamdaA => P(4)(218),lamdaB => P(4)(250),lamdaOut => P(3)(218));
F4219: entity F port map(lamdaA => P(4)(219),lamdaB => P(4)(251),lamdaOut => P(3)(219));
F4220: entity F port map(lamdaA => P(4)(220),lamdaB => P(4)(252),lamdaOut => P(3)(220));
F4221: entity F port map(lamdaA => P(4)(221),lamdaB => P(4)(253),lamdaOut => P(3)(221));
F4222: entity F port map(lamdaA => P(4)(222),lamdaB => P(4)(254),lamdaOut => P(3)(222));
F4223: entity F port map(lamdaA => P(4)(223),lamdaB => P(4)(255),lamdaOut => P(3)(223));
G4224: entity G port map(lamdaA => P(4)(192),lamdaB => P(4)(224),s => s(4)(96),lamdaOut => P(3)(224));
G4225: entity G port map(lamdaA => P(4)(193),lamdaB => P(4)(225),s => s(4)(97),lamdaOut => P(3)(225));
G4226: entity G port map(lamdaA => P(4)(194),lamdaB => P(4)(226),s => s(4)(98),lamdaOut => P(3)(226));
G4227: entity G port map(lamdaA => P(4)(195),lamdaB => P(4)(227),s => s(4)(99),lamdaOut => P(3)(227));
G4228: entity G port map(lamdaA => P(4)(196),lamdaB => P(4)(228),s => s(4)(100),lamdaOut => P(3)(228));
G4229: entity G port map(lamdaA => P(4)(197),lamdaB => P(4)(229),s => s(4)(101),lamdaOut => P(3)(229));
G4230: entity G port map(lamdaA => P(4)(198),lamdaB => P(4)(230),s => s(4)(102),lamdaOut => P(3)(230));
G4231: entity G port map(lamdaA => P(4)(199),lamdaB => P(4)(231),s => s(4)(103),lamdaOut => P(3)(231));
G4232: entity G port map(lamdaA => P(4)(200),lamdaB => P(4)(232),s => s(4)(104),lamdaOut => P(3)(232));
G4233: entity G port map(lamdaA => P(4)(201),lamdaB => P(4)(233),s => s(4)(105),lamdaOut => P(3)(233));
G4234: entity G port map(lamdaA => P(4)(202),lamdaB => P(4)(234),s => s(4)(106),lamdaOut => P(3)(234));
G4235: entity G port map(lamdaA => P(4)(203),lamdaB => P(4)(235),s => s(4)(107),lamdaOut => P(3)(235));
G4236: entity G port map(lamdaA => P(4)(204),lamdaB => P(4)(236),s => s(4)(108),lamdaOut => P(3)(236));
G4237: entity G port map(lamdaA => P(4)(205),lamdaB => P(4)(237),s => s(4)(109),lamdaOut => P(3)(237));
G4238: entity G port map(lamdaA => P(4)(206),lamdaB => P(4)(238),s => s(4)(110),lamdaOut => P(3)(238));
G4239: entity G port map(lamdaA => P(4)(207),lamdaB => P(4)(239),s => s(4)(111),lamdaOut => P(3)(239));
G4240: entity G port map(lamdaA => P(4)(208),lamdaB => P(4)(240),s => s(4)(112),lamdaOut => P(3)(240));
G4241: entity G port map(lamdaA => P(4)(209),lamdaB => P(4)(241),s => s(4)(113),lamdaOut => P(3)(241));
G4242: entity G port map(lamdaA => P(4)(210),lamdaB => P(4)(242),s => s(4)(114),lamdaOut => P(3)(242));
G4243: entity G port map(lamdaA => P(4)(211),lamdaB => P(4)(243),s => s(4)(115),lamdaOut => P(3)(243));
G4244: entity G port map(lamdaA => P(4)(212),lamdaB => P(4)(244),s => s(4)(116),lamdaOut => P(3)(244));
G4245: entity G port map(lamdaA => P(4)(213),lamdaB => P(4)(245),s => s(4)(117),lamdaOut => P(3)(245));
G4246: entity G port map(lamdaA => P(4)(214),lamdaB => P(4)(246),s => s(4)(118),lamdaOut => P(3)(246));
G4247: entity G port map(lamdaA => P(4)(215),lamdaB => P(4)(247),s => s(4)(119),lamdaOut => P(3)(247));
G4248: entity G port map(lamdaA => P(4)(216),lamdaB => P(4)(248),s => s(4)(120),lamdaOut => P(3)(248));
G4249: entity G port map(lamdaA => P(4)(217),lamdaB => P(4)(249),s => s(4)(121),lamdaOut => P(3)(249));
G4250: entity G port map(lamdaA => P(4)(218),lamdaB => P(4)(250),s => s(4)(122),lamdaOut => P(3)(250));
G4251: entity G port map(lamdaA => P(4)(219),lamdaB => P(4)(251),s => s(4)(123),lamdaOut => P(3)(251));
G4252: entity G port map(lamdaA => P(4)(220),lamdaB => P(4)(252),s => s(4)(124),lamdaOut => P(3)(252));
G4253: entity G port map(lamdaA => P(4)(221),lamdaB => P(4)(253),s => s(4)(125),lamdaOut => P(3)(253));
G4254: entity G port map(lamdaA => P(4)(222),lamdaB => P(4)(254),s => s(4)(126),lamdaOut => P(3)(254));
G4255: entity G port map(lamdaA => P(4)(223),lamdaB => P(4)(255),s => s(4)(127),lamdaOut => P(3)(255));
F4256: entity F port map(lamdaA => P(4)(256),lamdaB => P(4)(288),lamdaOut => P(3)(256));
F4257: entity F port map(lamdaA => P(4)(257),lamdaB => P(4)(289),lamdaOut => P(3)(257));
F4258: entity F port map(lamdaA => P(4)(258),lamdaB => P(4)(290),lamdaOut => P(3)(258));
F4259: entity F port map(lamdaA => P(4)(259),lamdaB => P(4)(291),lamdaOut => P(3)(259));
F4260: entity F port map(lamdaA => P(4)(260),lamdaB => P(4)(292),lamdaOut => P(3)(260));
F4261: entity F port map(lamdaA => P(4)(261),lamdaB => P(4)(293),lamdaOut => P(3)(261));
F4262: entity F port map(lamdaA => P(4)(262),lamdaB => P(4)(294),lamdaOut => P(3)(262));
F4263: entity F port map(lamdaA => P(4)(263),lamdaB => P(4)(295),lamdaOut => P(3)(263));
F4264: entity F port map(lamdaA => P(4)(264),lamdaB => P(4)(296),lamdaOut => P(3)(264));
F4265: entity F port map(lamdaA => P(4)(265),lamdaB => P(4)(297),lamdaOut => P(3)(265));
F4266: entity F port map(lamdaA => P(4)(266),lamdaB => P(4)(298),lamdaOut => P(3)(266));
F4267: entity F port map(lamdaA => P(4)(267),lamdaB => P(4)(299),lamdaOut => P(3)(267));
F4268: entity F port map(lamdaA => P(4)(268),lamdaB => P(4)(300),lamdaOut => P(3)(268));
F4269: entity F port map(lamdaA => P(4)(269),lamdaB => P(4)(301),lamdaOut => P(3)(269));
F4270: entity F port map(lamdaA => P(4)(270),lamdaB => P(4)(302),lamdaOut => P(3)(270));
F4271: entity F port map(lamdaA => P(4)(271),lamdaB => P(4)(303),lamdaOut => P(3)(271));
F4272: entity F port map(lamdaA => P(4)(272),lamdaB => P(4)(304),lamdaOut => P(3)(272));
F4273: entity F port map(lamdaA => P(4)(273),lamdaB => P(4)(305),lamdaOut => P(3)(273));
F4274: entity F port map(lamdaA => P(4)(274),lamdaB => P(4)(306),lamdaOut => P(3)(274));
F4275: entity F port map(lamdaA => P(4)(275),lamdaB => P(4)(307),lamdaOut => P(3)(275));
F4276: entity F port map(lamdaA => P(4)(276),lamdaB => P(4)(308),lamdaOut => P(3)(276));
F4277: entity F port map(lamdaA => P(4)(277),lamdaB => P(4)(309),lamdaOut => P(3)(277));
F4278: entity F port map(lamdaA => P(4)(278),lamdaB => P(4)(310),lamdaOut => P(3)(278));
F4279: entity F port map(lamdaA => P(4)(279),lamdaB => P(4)(311),lamdaOut => P(3)(279));
F4280: entity F port map(lamdaA => P(4)(280),lamdaB => P(4)(312),lamdaOut => P(3)(280));
F4281: entity F port map(lamdaA => P(4)(281),lamdaB => P(4)(313),lamdaOut => P(3)(281));
F4282: entity F port map(lamdaA => P(4)(282),lamdaB => P(4)(314),lamdaOut => P(3)(282));
F4283: entity F port map(lamdaA => P(4)(283),lamdaB => P(4)(315),lamdaOut => P(3)(283));
F4284: entity F port map(lamdaA => P(4)(284),lamdaB => P(4)(316),lamdaOut => P(3)(284));
F4285: entity F port map(lamdaA => P(4)(285),lamdaB => P(4)(317),lamdaOut => P(3)(285));
F4286: entity F port map(lamdaA => P(4)(286),lamdaB => P(4)(318),lamdaOut => P(3)(286));
F4287: entity F port map(lamdaA => P(4)(287),lamdaB => P(4)(319),lamdaOut => P(3)(287));
G4288: entity G port map(lamdaA => P(4)(256),lamdaB => P(4)(288),s => s(4)(128),lamdaOut => P(3)(288));
G4289: entity G port map(lamdaA => P(4)(257),lamdaB => P(4)(289),s => s(4)(129),lamdaOut => P(3)(289));
G4290: entity G port map(lamdaA => P(4)(258),lamdaB => P(4)(290),s => s(4)(130),lamdaOut => P(3)(290));
G4291: entity G port map(lamdaA => P(4)(259),lamdaB => P(4)(291),s => s(4)(131),lamdaOut => P(3)(291));
G4292: entity G port map(lamdaA => P(4)(260),lamdaB => P(4)(292),s => s(4)(132),lamdaOut => P(3)(292));
G4293: entity G port map(lamdaA => P(4)(261),lamdaB => P(4)(293),s => s(4)(133),lamdaOut => P(3)(293));
G4294: entity G port map(lamdaA => P(4)(262),lamdaB => P(4)(294),s => s(4)(134),lamdaOut => P(3)(294));
G4295: entity G port map(lamdaA => P(4)(263),lamdaB => P(4)(295),s => s(4)(135),lamdaOut => P(3)(295));
G4296: entity G port map(lamdaA => P(4)(264),lamdaB => P(4)(296),s => s(4)(136),lamdaOut => P(3)(296));
G4297: entity G port map(lamdaA => P(4)(265),lamdaB => P(4)(297),s => s(4)(137),lamdaOut => P(3)(297));
G4298: entity G port map(lamdaA => P(4)(266),lamdaB => P(4)(298),s => s(4)(138),lamdaOut => P(3)(298));
G4299: entity G port map(lamdaA => P(4)(267),lamdaB => P(4)(299),s => s(4)(139),lamdaOut => P(3)(299));
G4300: entity G port map(lamdaA => P(4)(268),lamdaB => P(4)(300),s => s(4)(140),lamdaOut => P(3)(300));
G4301: entity G port map(lamdaA => P(4)(269),lamdaB => P(4)(301),s => s(4)(141),lamdaOut => P(3)(301));
G4302: entity G port map(lamdaA => P(4)(270),lamdaB => P(4)(302),s => s(4)(142),lamdaOut => P(3)(302));
G4303: entity G port map(lamdaA => P(4)(271),lamdaB => P(4)(303),s => s(4)(143),lamdaOut => P(3)(303));
G4304: entity G port map(lamdaA => P(4)(272),lamdaB => P(4)(304),s => s(4)(144),lamdaOut => P(3)(304));
G4305: entity G port map(lamdaA => P(4)(273),lamdaB => P(4)(305),s => s(4)(145),lamdaOut => P(3)(305));
G4306: entity G port map(lamdaA => P(4)(274),lamdaB => P(4)(306),s => s(4)(146),lamdaOut => P(3)(306));
G4307: entity G port map(lamdaA => P(4)(275),lamdaB => P(4)(307),s => s(4)(147),lamdaOut => P(3)(307));
G4308: entity G port map(lamdaA => P(4)(276),lamdaB => P(4)(308),s => s(4)(148),lamdaOut => P(3)(308));
G4309: entity G port map(lamdaA => P(4)(277),lamdaB => P(4)(309),s => s(4)(149),lamdaOut => P(3)(309));
G4310: entity G port map(lamdaA => P(4)(278),lamdaB => P(4)(310),s => s(4)(150),lamdaOut => P(3)(310));
G4311: entity G port map(lamdaA => P(4)(279),lamdaB => P(4)(311),s => s(4)(151),lamdaOut => P(3)(311));
G4312: entity G port map(lamdaA => P(4)(280),lamdaB => P(4)(312),s => s(4)(152),lamdaOut => P(3)(312));
G4313: entity G port map(lamdaA => P(4)(281),lamdaB => P(4)(313),s => s(4)(153),lamdaOut => P(3)(313));
G4314: entity G port map(lamdaA => P(4)(282),lamdaB => P(4)(314),s => s(4)(154),lamdaOut => P(3)(314));
G4315: entity G port map(lamdaA => P(4)(283),lamdaB => P(4)(315),s => s(4)(155),lamdaOut => P(3)(315));
G4316: entity G port map(lamdaA => P(4)(284),lamdaB => P(4)(316),s => s(4)(156),lamdaOut => P(3)(316));
G4317: entity G port map(lamdaA => P(4)(285),lamdaB => P(4)(317),s => s(4)(157),lamdaOut => P(3)(317));
G4318: entity G port map(lamdaA => P(4)(286),lamdaB => P(4)(318),s => s(4)(158),lamdaOut => P(3)(318));
G4319: entity G port map(lamdaA => P(4)(287),lamdaB => P(4)(319),s => s(4)(159),lamdaOut => P(3)(319));
F4320: entity F port map(lamdaA => P(4)(320),lamdaB => P(4)(352),lamdaOut => P(3)(320));
F4321: entity F port map(lamdaA => P(4)(321),lamdaB => P(4)(353),lamdaOut => P(3)(321));
F4322: entity F port map(lamdaA => P(4)(322),lamdaB => P(4)(354),lamdaOut => P(3)(322));
F4323: entity F port map(lamdaA => P(4)(323),lamdaB => P(4)(355),lamdaOut => P(3)(323));
F4324: entity F port map(lamdaA => P(4)(324),lamdaB => P(4)(356),lamdaOut => P(3)(324));
F4325: entity F port map(lamdaA => P(4)(325),lamdaB => P(4)(357),lamdaOut => P(3)(325));
F4326: entity F port map(lamdaA => P(4)(326),lamdaB => P(4)(358),lamdaOut => P(3)(326));
F4327: entity F port map(lamdaA => P(4)(327),lamdaB => P(4)(359),lamdaOut => P(3)(327));
F4328: entity F port map(lamdaA => P(4)(328),lamdaB => P(4)(360),lamdaOut => P(3)(328));
F4329: entity F port map(lamdaA => P(4)(329),lamdaB => P(4)(361),lamdaOut => P(3)(329));
F4330: entity F port map(lamdaA => P(4)(330),lamdaB => P(4)(362),lamdaOut => P(3)(330));
F4331: entity F port map(lamdaA => P(4)(331),lamdaB => P(4)(363),lamdaOut => P(3)(331));
F4332: entity F port map(lamdaA => P(4)(332),lamdaB => P(4)(364),lamdaOut => P(3)(332));
F4333: entity F port map(lamdaA => P(4)(333),lamdaB => P(4)(365),lamdaOut => P(3)(333));
F4334: entity F port map(lamdaA => P(4)(334),lamdaB => P(4)(366),lamdaOut => P(3)(334));
F4335: entity F port map(lamdaA => P(4)(335),lamdaB => P(4)(367),lamdaOut => P(3)(335));
F4336: entity F port map(lamdaA => P(4)(336),lamdaB => P(4)(368),lamdaOut => P(3)(336));
F4337: entity F port map(lamdaA => P(4)(337),lamdaB => P(4)(369),lamdaOut => P(3)(337));
F4338: entity F port map(lamdaA => P(4)(338),lamdaB => P(4)(370),lamdaOut => P(3)(338));
F4339: entity F port map(lamdaA => P(4)(339),lamdaB => P(4)(371),lamdaOut => P(3)(339));
F4340: entity F port map(lamdaA => P(4)(340),lamdaB => P(4)(372),lamdaOut => P(3)(340));
F4341: entity F port map(lamdaA => P(4)(341),lamdaB => P(4)(373),lamdaOut => P(3)(341));
F4342: entity F port map(lamdaA => P(4)(342),lamdaB => P(4)(374),lamdaOut => P(3)(342));
F4343: entity F port map(lamdaA => P(4)(343),lamdaB => P(4)(375),lamdaOut => P(3)(343));
F4344: entity F port map(lamdaA => P(4)(344),lamdaB => P(4)(376),lamdaOut => P(3)(344));
F4345: entity F port map(lamdaA => P(4)(345),lamdaB => P(4)(377),lamdaOut => P(3)(345));
F4346: entity F port map(lamdaA => P(4)(346),lamdaB => P(4)(378),lamdaOut => P(3)(346));
F4347: entity F port map(lamdaA => P(4)(347),lamdaB => P(4)(379),lamdaOut => P(3)(347));
F4348: entity F port map(lamdaA => P(4)(348),lamdaB => P(4)(380),lamdaOut => P(3)(348));
F4349: entity F port map(lamdaA => P(4)(349),lamdaB => P(4)(381),lamdaOut => P(3)(349));
F4350: entity F port map(lamdaA => P(4)(350),lamdaB => P(4)(382),lamdaOut => P(3)(350));
F4351: entity F port map(lamdaA => P(4)(351),lamdaB => P(4)(383),lamdaOut => P(3)(351));
G4352: entity G port map(lamdaA => P(4)(320),lamdaB => P(4)(352),s => s(4)(160),lamdaOut => P(3)(352));
G4353: entity G port map(lamdaA => P(4)(321),lamdaB => P(4)(353),s => s(4)(161),lamdaOut => P(3)(353));
G4354: entity G port map(lamdaA => P(4)(322),lamdaB => P(4)(354),s => s(4)(162),lamdaOut => P(3)(354));
G4355: entity G port map(lamdaA => P(4)(323),lamdaB => P(4)(355),s => s(4)(163),lamdaOut => P(3)(355));
G4356: entity G port map(lamdaA => P(4)(324),lamdaB => P(4)(356),s => s(4)(164),lamdaOut => P(3)(356));
G4357: entity G port map(lamdaA => P(4)(325),lamdaB => P(4)(357),s => s(4)(165),lamdaOut => P(3)(357));
G4358: entity G port map(lamdaA => P(4)(326),lamdaB => P(4)(358),s => s(4)(166),lamdaOut => P(3)(358));
G4359: entity G port map(lamdaA => P(4)(327),lamdaB => P(4)(359),s => s(4)(167),lamdaOut => P(3)(359));
G4360: entity G port map(lamdaA => P(4)(328),lamdaB => P(4)(360),s => s(4)(168),lamdaOut => P(3)(360));
G4361: entity G port map(lamdaA => P(4)(329),lamdaB => P(4)(361),s => s(4)(169),lamdaOut => P(3)(361));
G4362: entity G port map(lamdaA => P(4)(330),lamdaB => P(4)(362),s => s(4)(170),lamdaOut => P(3)(362));
G4363: entity G port map(lamdaA => P(4)(331),lamdaB => P(4)(363),s => s(4)(171),lamdaOut => P(3)(363));
G4364: entity G port map(lamdaA => P(4)(332),lamdaB => P(4)(364),s => s(4)(172),lamdaOut => P(3)(364));
G4365: entity G port map(lamdaA => P(4)(333),lamdaB => P(4)(365),s => s(4)(173),lamdaOut => P(3)(365));
G4366: entity G port map(lamdaA => P(4)(334),lamdaB => P(4)(366),s => s(4)(174),lamdaOut => P(3)(366));
G4367: entity G port map(lamdaA => P(4)(335),lamdaB => P(4)(367),s => s(4)(175),lamdaOut => P(3)(367));
G4368: entity G port map(lamdaA => P(4)(336),lamdaB => P(4)(368),s => s(4)(176),lamdaOut => P(3)(368));
G4369: entity G port map(lamdaA => P(4)(337),lamdaB => P(4)(369),s => s(4)(177),lamdaOut => P(3)(369));
G4370: entity G port map(lamdaA => P(4)(338),lamdaB => P(4)(370),s => s(4)(178),lamdaOut => P(3)(370));
G4371: entity G port map(lamdaA => P(4)(339),lamdaB => P(4)(371),s => s(4)(179),lamdaOut => P(3)(371));
G4372: entity G port map(lamdaA => P(4)(340),lamdaB => P(4)(372),s => s(4)(180),lamdaOut => P(3)(372));
G4373: entity G port map(lamdaA => P(4)(341),lamdaB => P(4)(373),s => s(4)(181),lamdaOut => P(3)(373));
G4374: entity G port map(lamdaA => P(4)(342),lamdaB => P(4)(374),s => s(4)(182),lamdaOut => P(3)(374));
G4375: entity G port map(lamdaA => P(4)(343),lamdaB => P(4)(375),s => s(4)(183),lamdaOut => P(3)(375));
G4376: entity G port map(lamdaA => P(4)(344),lamdaB => P(4)(376),s => s(4)(184),lamdaOut => P(3)(376));
G4377: entity G port map(lamdaA => P(4)(345),lamdaB => P(4)(377),s => s(4)(185),lamdaOut => P(3)(377));
G4378: entity G port map(lamdaA => P(4)(346),lamdaB => P(4)(378),s => s(4)(186),lamdaOut => P(3)(378));
G4379: entity G port map(lamdaA => P(4)(347),lamdaB => P(4)(379),s => s(4)(187),lamdaOut => P(3)(379));
G4380: entity G port map(lamdaA => P(4)(348),lamdaB => P(4)(380),s => s(4)(188),lamdaOut => P(3)(380));
G4381: entity G port map(lamdaA => P(4)(349),lamdaB => P(4)(381),s => s(4)(189),lamdaOut => P(3)(381));
G4382: entity G port map(lamdaA => P(4)(350),lamdaB => P(4)(382),s => s(4)(190),lamdaOut => P(3)(382));
G4383: entity G port map(lamdaA => P(4)(351),lamdaB => P(4)(383),s => s(4)(191),lamdaOut => P(3)(383));
F4384: entity F port map(lamdaA => P(4)(384),lamdaB => P(4)(416),lamdaOut => P(3)(384));
F4385: entity F port map(lamdaA => P(4)(385),lamdaB => P(4)(417),lamdaOut => P(3)(385));
F4386: entity F port map(lamdaA => P(4)(386),lamdaB => P(4)(418),lamdaOut => P(3)(386));
F4387: entity F port map(lamdaA => P(4)(387),lamdaB => P(4)(419),lamdaOut => P(3)(387));
F4388: entity F port map(lamdaA => P(4)(388),lamdaB => P(4)(420),lamdaOut => P(3)(388));
F4389: entity F port map(lamdaA => P(4)(389),lamdaB => P(4)(421),lamdaOut => P(3)(389));
F4390: entity F port map(lamdaA => P(4)(390),lamdaB => P(4)(422),lamdaOut => P(3)(390));
F4391: entity F port map(lamdaA => P(4)(391),lamdaB => P(4)(423),lamdaOut => P(3)(391));
F4392: entity F port map(lamdaA => P(4)(392),lamdaB => P(4)(424),lamdaOut => P(3)(392));
F4393: entity F port map(lamdaA => P(4)(393),lamdaB => P(4)(425),lamdaOut => P(3)(393));
F4394: entity F port map(lamdaA => P(4)(394),lamdaB => P(4)(426),lamdaOut => P(3)(394));
F4395: entity F port map(lamdaA => P(4)(395),lamdaB => P(4)(427),lamdaOut => P(3)(395));
F4396: entity F port map(lamdaA => P(4)(396),lamdaB => P(4)(428),lamdaOut => P(3)(396));
F4397: entity F port map(lamdaA => P(4)(397),lamdaB => P(4)(429),lamdaOut => P(3)(397));
F4398: entity F port map(lamdaA => P(4)(398),lamdaB => P(4)(430),lamdaOut => P(3)(398));
F4399: entity F port map(lamdaA => P(4)(399),lamdaB => P(4)(431),lamdaOut => P(3)(399));
F4400: entity F port map(lamdaA => P(4)(400),lamdaB => P(4)(432),lamdaOut => P(3)(400));
F4401: entity F port map(lamdaA => P(4)(401),lamdaB => P(4)(433),lamdaOut => P(3)(401));
F4402: entity F port map(lamdaA => P(4)(402),lamdaB => P(4)(434),lamdaOut => P(3)(402));
F4403: entity F port map(lamdaA => P(4)(403),lamdaB => P(4)(435),lamdaOut => P(3)(403));
F4404: entity F port map(lamdaA => P(4)(404),lamdaB => P(4)(436),lamdaOut => P(3)(404));
F4405: entity F port map(lamdaA => P(4)(405),lamdaB => P(4)(437),lamdaOut => P(3)(405));
F4406: entity F port map(lamdaA => P(4)(406),lamdaB => P(4)(438),lamdaOut => P(3)(406));
F4407: entity F port map(lamdaA => P(4)(407),lamdaB => P(4)(439),lamdaOut => P(3)(407));
F4408: entity F port map(lamdaA => P(4)(408),lamdaB => P(4)(440),lamdaOut => P(3)(408));
F4409: entity F port map(lamdaA => P(4)(409),lamdaB => P(4)(441),lamdaOut => P(3)(409));
F4410: entity F port map(lamdaA => P(4)(410),lamdaB => P(4)(442),lamdaOut => P(3)(410));
F4411: entity F port map(lamdaA => P(4)(411),lamdaB => P(4)(443),lamdaOut => P(3)(411));
F4412: entity F port map(lamdaA => P(4)(412),lamdaB => P(4)(444),lamdaOut => P(3)(412));
F4413: entity F port map(lamdaA => P(4)(413),lamdaB => P(4)(445),lamdaOut => P(3)(413));
F4414: entity F port map(lamdaA => P(4)(414),lamdaB => P(4)(446),lamdaOut => P(3)(414));
F4415: entity F port map(lamdaA => P(4)(415),lamdaB => P(4)(447),lamdaOut => P(3)(415));
G4416: entity G port map(lamdaA => P(4)(384),lamdaB => P(4)(416),s => s(4)(192),lamdaOut => P(3)(416));
G4417: entity G port map(lamdaA => P(4)(385),lamdaB => P(4)(417),s => s(4)(193),lamdaOut => P(3)(417));
G4418: entity G port map(lamdaA => P(4)(386),lamdaB => P(4)(418),s => s(4)(194),lamdaOut => P(3)(418));
G4419: entity G port map(lamdaA => P(4)(387),lamdaB => P(4)(419),s => s(4)(195),lamdaOut => P(3)(419));
G4420: entity G port map(lamdaA => P(4)(388),lamdaB => P(4)(420),s => s(4)(196),lamdaOut => P(3)(420));
G4421: entity G port map(lamdaA => P(4)(389),lamdaB => P(4)(421),s => s(4)(197),lamdaOut => P(3)(421));
G4422: entity G port map(lamdaA => P(4)(390),lamdaB => P(4)(422),s => s(4)(198),lamdaOut => P(3)(422));
G4423: entity G port map(lamdaA => P(4)(391),lamdaB => P(4)(423),s => s(4)(199),lamdaOut => P(3)(423));
G4424: entity G port map(lamdaA => P(4)(392),lamdaB => P(4)(424),s => s(4)(200),lamdaOut => P(3)(424));
G4425: entity G port map(lamdaA => P(4)(393),lamdaB => P(4)(425),s => s(4)(201),lamdaOut => P(3)(425));
G4426: entity G port map(lamdaA => P(4)(394),lamdaB => P(4)(426),s => s(4)(202),lamdaOut => P(3)(426));
G4427: entity G port map(lamdaA => P(4)(395),lamdaB => P(4)(427),s => s(4)(203),lamdaOut => P(3)(427));
G4428: entity G port map(lamdaA => P(4)(396),lamdaB => P(4)(428),s => s(4)(204),lamdaOut => P(3)(428));
G4429: entity G port map(lamdaA => P(4)(397),lamdaB => P(4)(429),s => s(4)(205),lamdaOut => P(3)(429));
G4430: entity G port map(lamdaA => P(4)(398),lamdaB => P(4)(430),s => s(4)(206),lamdaOut => P(3)(430));
G4431: entity G port map(lamdaA => P(4)(399),lamdaB => P(4)(431),s => s(4)(207),lamdaOut => P(3)(431));
G4432: entity G port map(lamdaA => P(4)(400),lamdaB => P(4)(432),s => s(4)(208),lamdaOut => P(3)(432));
G4433: entity G port map(lamdaA => P(4)(401),lamdaB => P(4)(433),s => s(4)(209),lamdaOut => P(3)(433));
G4434: entity G port map(lamdaA => P(4)(402),lamdaB => P(4)(434),s => s(4)(210),lamdaOut => P(3)(434));
G4435: entity G port map(lamdaA => P(4)(403),lamdaB => P(4)(435),s => s(4)(211),lamdaOut => P(3)(435));
G4436: entity G port map(lamdaA => P(4)(404),lamdaB => P(4)(436),s => s(4)(212),lamdaOut => P(3)(436));
G4437: entity G port map(lamdaA => P(4)(405),lamdaB => P(4)(437),s => s(4)(213),lamdaOut => P(3)(437));
G4438: entity G port map(lamdaA => P(4)(406),lamdaB => P(4)(438),s => s(4)(214),lamdaOut => P(3)(438));
G4439: entity G port map(lamdaA => P(4)(407),lamdaB => P(4)(439),s => s(4)(215),lamdaOut => P(3)(439));
G4440: entity G port map(lamdaA => P(4)(408),lamdaB => P(4)(440),s => s(4)(216),lamdaOut => P(3)(440));
G4441: entity G port map(lamdaA => P(4)(409),lamdaB => P(4)(441),s => s(4)(217),lamdaOut => P(3)(441));
G4442: entity G port map(lamdaA => P(4)(410),lamdaB => P(4)(442),s => s(4)(218),lamdaOut => P(3)(442));
G4443: entity G port map(lamdaA => P(4)(411),lamdaB => P(4)(443),s => s(4)(219),lamdaOut => P(3)(443));
G4444: entity G port map(lamdaA => P(4)(412),lamdaB => P(4)(444),s => s(4)(220),lamdaOut => P(3)(444));
G4445: entity G port map(lamdaA => P(4)(413),lamdaB => P(4)(445),s => s(4)(221),lamdaOut => P(3)(445));
G4446: entity G port map(lamdaA => P(4)(414),lamdaB => P(4)(446),s => s(4)(222),lamdaOut => P(3)(446));
G4447: entity G port map(lamdaA => P(4)(415),lamdaB => P(4)(447),s => s(4)(223),lamdaOut => P(3)(447));
F4448: entity F port map(lamdaA => P(4)(448),lamdaB => P(4)(480),lamdaOut => P(3)(448));
F4449: entity F port map(lamdaA => P(4)(449),lamdaB => P(4)(481),lamdaOut => P(3)(449));
F4450: entity F port map(lamdaA => P(4)(450),lamdaB => P(4)(482),lamdaOut => P(3)(450));
F4451: entity F port map(lamdaA => P(4)(451),lamdaB => P(4)(483),lamdaOut => P(3)(451));
F4452: entity F port map(lamdaA => P(4)(452),lamdaB => P(4)(484),lamdaOut => P(3)(452));
F4453: entity F port map(lamdaA => P(4)(453),lamdaB => P(4)(485),lamdaOut => P(3)(453));
F4454: entity F port map(lamdaA => P(4)(454),lamdaB => P(4)(486),lamdaOut => P(3)(454));
F4455: entity F port map(lamdaA => P(4)(455),lamdaB => P(4)(487),lamdaOut => P(3)(455));
F4456: entity F port map(lamdaA => P(4)(456),lamdaB => P(4)(488),lamdaOut => P(3)(456));
F4457: entity F port map(lamdaA => P(4)(457),lamdaB => P(4)(489),lamdaOut => P(3)(457));
F4458: entity F port map(lamdaA => P(4)(458),lamdaB => P(4)(490),lamdaOut => P(3)(458));
F4459: entity F port map(lamdaA => P(4)(459),lamdaB => P(4)(491),lamdaOut => P(3)(459));
F4460: entity F port map(lamdaA => P(4)(460),lamdaB => P(4)(492),lamdaOut => P(3)(460));
F4461: entity F port map(lamdaA => P(4)(461),lamdaB => P(4)(493),lamdaOut => P(3)(461));
F4462: entity F port map(lamdaA => P(4)(462),lamdaB => P(4)(494),lamdaOut => P(3)(462));
F4463: entity F port map(lamdaA => P(4)(463),lamdaB => P(4)(495),lamdaOut => P(3)(463));
F4464: entity F port map(lamdaA => P(4)(464),lamdaB => P(4)(496),lamdaOut => P(3)(464));
F4465: entity F port map(lamdaA => P(4)(465),lamdaB => P(4)(497),lamdaOut => P(3)(465));
F4466: entity F port map(lamdaA => P(4)(466),lamdaB => P(4)(498),lamdaOut => P(3)(466));
F4467: entity F port map(lamdaA => P(4)(467),lamdaB => P(4)(499),lamdaOut => P(3)(467));
F4468: entity F port map(lamdaA => P(4)(468),lamdaB => P(4)(500),lamdaOut => P(3)(468));
F4469: entity F port map(lamdaA => P(4)(469),lamdaB => P(4)(501),lamdaOut => P(3)(469));
F4470: entity F port map(lamdaA => P(4)(470),lamdaB => P(4)(502),lamdaOut => P(3)(470));
F4471: entity F port map(lamdaA => P(4)(471),lamdaB => P(4)(503),lamdaOut => P(3)(471));
F4472: entity F port map(lamdaA => P(4)(472),lamdaB => P(4)(504),lamdaOut => P(3)(472));
F4473: entity F port map(lamdaA => P(4)(473),lamdaB => P(4)(505),lamdaOut => P(3)(473));
F4474: entity F port map(lamdaA => P(4)(474),lamdaB => P(4)(506),lamdaOut => P(3)(474));
F4475: entity F port map(lamdaA => P(4)(475),lamdaB => P(4)(507),lamdaOut => P(3)(475));
F4476: entity F port map(lamdaA => P(4)(476),lamdaB => P(4)(508),lamdaOut => P(3)(476));
F4477: entity F port map(lamdaA => P(4)(477),lamdaB => P(4)(509),lamdaOut => P(3)(477));
F4478: entity F port map(lamdaA => P(4)(478),lamdaB => P(4)(510),lamdaOut => P(3)(478));
F4479: entity F port map(lamdaA => P(4)(479),lamdaB => P(4)(511),lamdaOut => P(3)(479));
G4480: entity G port map(lamdaA => P(4)(448),lamdaB => P(4)(480),s => s(4)(224),lamdaOut => P(3)(480));
G4481: entity G port map(lamdaA => P(4)(449),lamdaB => P(4)(481),s => s(4)(225),lamdaOut => P(3)(481));
G4482: entity G port map(lamdaA => P(4)(450),lamdaB => P(4)(482),s => s(4)(226),lamdaOut => P(3)(482));
G4483: entity G port map(lamdaA => P(4)(451),lamdaB => P(4)(483),s => s(4)(227),lamdaOut => P(3)(483));
G4484: entity G port map(lamdaA => P(4)(452),lamdaB => P(4)(484),s => s(4)(228),lamdaOut => P(3)(484));
G4485: entity G port map(lamdaA => P(4)(453),lamdaB => P(4)(485),s => s(4)(229),lamdaOut => P(3)(485));
G4486: entity G port map(lamdaA => P(4)(454),lamdaB => P(4)(486),s => s(4)(230),lamdaOut => P(3)(486));
G4487: entity G port map(lamdaA => P(4)(455),lamdaB => P(4)(487),s => s(4)(231),lamdaOut => P(3)(487));
G4488: entity G port map(lamdaA => P(4)(456),lamdaB => P(4)(488),s => s(4)(232),lamdaOut => P(3)(488));
G4489: entity G port map(lamdaA => P(4)(457),lamdaB => P(4)(489),s => s(4)(233),lamdaOut => P(3)(489));
G4490: entity G port map(lamdaA => P(4)(458),lamdaB => P(4)(490),s => s(4)(234),lamdaOut => P(3)(490));
G4491: entity G port map(lamdaA => P(4)(459),lamdaB => P(4)(491),s => s(4)(235),lamdaOut => P(3)(491));
G4492: entity G port map(lamdaA => P(4)(460),lamdaB => P(4)(492),s => s(4)(236),lamdaOut => P(3)(492));
G4493: entity G port map(lamdaA => P(4)(461),lamdaB => P(4)(493),s => s(4)(237),lamdaOut => P(3)(493));
G4494: entity G port map(lamdaA => P(4)(462),lamdaB => P(4)(494),s => s(4)(238),lamdaOut => P(3)(494));
G4495: entity G port map(lamdaA => P(4)(463),lamdaB => P(4)(495),s => s(4)(239),lamdaOut => P(3)(495));
G4496: entity G port map(lamdaA => P(4)(464),lamdaB => P(4)(496),s => s(4)(240),lamdaOut => P(3)(496));
G4497: entity G port map(lamdaA => P(4)(465),lamdaB => P(4)(497),s => s(4)(241),lamdaOut => P(3)(497));
G4498: entity G port map(lamdaA => P(4)(466),lamdaB => P(4)(498),s => s(4)(242),lamdaOut => P(3)(498));
G4499: entity G port map(lamdaA => P(4)(467),lamdaB => P(4)(499),s => s(4)(243),lamdaOut => P(3)(499));
G4500: entity G port map(lamdaA => P(4)(468),lamdaB => P(4)(500),s => s(4)(244),lamdaOut => P(3)(500));
G4501: entity G port map(lamdaA => P(4)(469),lamdaB => P(4)(501),s => s(4)(245),lamdaOut => P(3)(501));
G4502: entity G port map(lamdaA => P(4)(470),lamdaB => P(4)(502),s => s(4)(246),lamdaOut => P(3)(502));
G4503: entity G port map(lamdaA => P(4)(471),lamdaB => P(4)(503),s => s(4)(247),lamdaOut => P(3)(503));
G4504: entity G port map(lamdaA => P(4)(472),lamdaB => P(4)(504),s => s(4)(248),lamdaOut => P(3)(504));
G4505: entity G port map(lamdaA => P(4)(473),lamdaB => P(4)(505),s => s(4)(249),lamdaOut => P(3)(505));
G4506: entity G port map(lamdaA => P(4)(474),lamdaB => P(4)(506),s => s(4)(250),lamdaOut => P(3)(506));
G4507: entity G port map(lamdaA => P(4)(475),lamdaB => P(4)(507),s => s(4)(251),lamdaOut => P(3)(507));
G4508: entity G port map(lamdaA => P(4)(476),lamdaB => P(4)(508),s => s(4)(252),lamdaOut => P(3)(508));
G4509: entity G port map(lamdaA => P(4)(477),lamdaB => P(4)(509),s => s(4)(253),lamdaOut => P(3)(509));
G4510: entity G port map(lamdaA => P(4)(478),lamdaB => P(4)(510),s => s(4)(254),lamdaOut => P(3)(510));
G4511: entity G port map(lamdaA => P(4)(479),lamdaB => P(4)(511),s => s(4)(255),lamdaOut => P(3)(511));
-- STAGE 3
F30: entity F port map(lamdaA => P(3)(0),lamdaB => P(3)(64),lamdaOut => P(2)(0));
F31: entity F port map(lamdaA => P(3)(1),lamdaB => P(3)(65),lamdaOut => P(2)(1));
F32: entity F port map(lamdaA => P(3)(2),lamdaB => P(3)(66),lamdaOut => P(2)(2));
F33: entity F port map(lamdaA => P(3)(3),lamdaB => P(3)(67),lamdaOut => P(2)(3));
F34: entity F port map(lamdaA => P(3)(4),lamdaB => P(3)(68),lamdaOut => P(2)(4));
F35: entity F port map(lamdaA => P(3)(5),lamdaB => P(3)(69),lamdaOut => P(2)(5));
F36: entity F port map(lamdaA => P(3)(6),lamdaB => P(3)(70),lamdaOut => P(2)(6));
F37: entity F port map(lamdaA => P(3)(7),lamdaB => P(3)(71),lamdaOut => P(2)(7));
F38: entity F port map(lamdaA => P(3)(8),lamdaB => P(3)(72),lamdaOut => P(2)(8));
F39: entity F port map(lamdaA => P(3)(9),lamdaB => P(3)(73),lamdaOut => P(2)(9));
F310: entity F port map(lamdaA => P(3)(10),lamdaB => P(3)(74),lamdaOut => P(2)(10));
F311: entity F port map(lamdaA => P(3)(11),lamdaB => P(3)(75),lamdaOut => P(2)(11));
F312: entity F port map(lamdaA => P(3)(12),lamdaB => P(3)(76),lamdaOut => P(2)(12));
F313: entity F port map(lamdaA => P(3)(13),lamdaB => P(3)(77),lamdaOut => P(2)(13));
F314: entity F port map(lamdaA => P(3)(14),lamdaB => P(3)(78),lamdaOut => P(2)(14));
F315: entity F port map(lamdaA => P(3)(15),lamdaB => P(3)(79),lamdaOut => P(2)(15));
F316: entity F port map(lamdaA => P(3)(16),lamdaB => P(3)(80),lamdaOut => P(2)(16));
F317: entity F port map(lamdaA => P(3)(17),lamdaB => P(3)(81),lamdaOut => P(2)(17));
F318: entity F port map(lamdaA => P(3)(18),lamdaB => P(3)(82),lamdaOut => P(2)(18));
F319: entity F port map(lamdaA => P(3)(19),lamdaB => P(3)(83),lamdaOut => P(2)(19));
F320: entity F port map(lamdaA => P(3)(20),lamdaB => P(3)(84),lamdaOut => P(2)(20));
F321: entity F port map(lamdaA => P(3)(21),lamdaB => P(3)(85),lamdaOut => P(2)(21));
F322: entity F port map(lamdaA => P(3)(22),lamdaB => P(3)(86),lamdaOut => P(2)(22));
F323: entity F port map(lamdaA => P(3)(23),lamdaB => P(3)(87),lamdaOut => P(2)(23));
F324: entity F port map(lamdaA => P(3)(24),lamdaB => P(3)(88),lamdaOut => P(2)(24));
F325: entity F port map(lamdaA => P(3)(25),lamdaB => P(3)(89),lamdaOut => P(2)(25));
F326: entity F port map(lamdaA => P(3)(26),lamdaB => P(3)(90),lamdaOut => P(2)(26));
F327: entity F port map(lamdaA => P(3)(27),lamdaB => P(3)(91),lamdaOut => P(2)(27));
F328: entity F port map(lamdaA => P(3)(28),lamdaB => P(3)(92),lamdaOut => P(2)(28));
F329: entity F port map(lamdaA => P(3)(29),lamdaB => P(3)(93),lamdaOut => P(2)(29));
F330: entity F port map(lamdaA => P(3)(30),lamdaB => P(3)(94),lamdaOut => P(2)(30));
F331: entity F port map(lamdaA => P(3)(31),lamdaB => P(3)(95),lamdaOut => P(2)(31));
F332: entity F port map(lamdaA => P(3)(32),lamdaB => P(3)(96),lamdaOut => P(2)(32));
F333: entity F port map(lamdaA => P(3)(33),lamdaB => P(3)(97),lamdaOut => P(2)(33));
F334: entity F port map(lamdaA => P(3)(34),lamdaB => P(3)(98),lamdaOut => P(2)(34));
F335: entity F port map(lamdaA => P(3)(35),lamdaB => P(3)(99),lamdaOut => P(2)(35));
F336: entity F port map(lamdaA => P(3)(36),lamdaB => P(3)(100),lamdaOut => P(2)(36));
F337: entity F port map(lamdaA => P(3)(37),lamdaB => P(3)(101),lamdaOut => P(2)(37));
F338: entity F port map(lamdaA => P(3)(38),lamdaB => P(3)(102),lamdaOut => P(2)(38));
F339: entity F port map(lamdaA => P(3)(39),lamdaB => P(3)(103),lamdaOut => P(2)(39));
F340: entity F port map(lamdaA => P(3)(40),lamdaB => P(3)(104),lamdaOut => P(2)(40));
F341: entity F port map(lamdaA => P(3)(41),lamdaB => P(3)(105),lamdaOut => P(2)(41));
F342: entity F port map(lamdaA => P(3)(42),lamdaB => P(3)(106),lamdaOut => P(2)(42));
F343: entity F port map(lamdaA => P(3)(43),lamdaB => P(3)(107),lamdaOut => P(2)(43));
F344: entity F port map(lamdaA => P(3)(44),lamdaB => P(3)(108),lamdaOut => P(2)(44));
F345: entity F port map(lamdaA => P(3)(45),lamdaB => P(3)(109),lamdaOut => P(2)(45));
F346: entity F port map(lamdaA => P(3)(46),lamdaB => P(3)(110),lamdaOut => P(2)(46));
F347: entity F port map(lamdaA => P(3)(47),lamdaB => P(3)(111),lamdaOut => P(2)(47));
F348: entity F port map(lamdaA => P(3)(48),lamdaB => P(3)(112),lamdaOut => P(2)(48));
F349: entity F port map(lamdaA => P(3)(49),lamdaB => P(3)(113),lamdaOut => P(2)(49));
F350: entity F port map(lamdaA => P(3)(50),lamdaB => P(3)(114),lamdaOut => P(2)(50));
F351: entity F port map(lamdaA => P(3)(51),lamdaB => P(3)(115),lamdaOut => P(2)(51));
F352: entity F port map(lamdaA => P(3)(52),lamdaB => P(3)(116),lamdaOut => P(2)(52));
F353: entity F port map(lamdaA => P(3)(53),lamdaB => P(3)(117),lamdaOut => P(2)(53));
F354: entity F port map(lamdaA => P(3)(54),lamdaB => P(3)(118),lamdaOut => P(2)(54));
F355: entity F port map(lamdaA => P(3)(55),lamdaB => P(3)(119),lamdaOut => P(2)(55));
F356: entity F port map(lamdaA => P(3)(56),lamdaB => P(3)(120),lamdaOut => P(2)(56));
F357: entity F port map(lamdaA => P(3)(57),lamdaB => P(3)(121),lamdaOut => P(2)(57));
F358: entity F port map(lamdaA => P(3)(58),lamdaB => P(3)(122),lamdaOut => P(2)(58));
F359: entity F port map(lamdaA => P(3)(59),lamdaB => P(3)(123),lamdaOut => P(2)(59));
F360: entity F port map(lamdaA => P(3)(60),lamdaB => P(3)(124),lamdaOut => P(2)(60));
F361: entity F port map(lamdaA => P(3)(61),lamdaB => P(3)(125),lamdaOut => P(2)(61));
F362: entity F port map(lamdaA => P(3)(62),lamdaB => P(3)(126),lamdaOut => P(2)(62));
F363: entity F port map(lamdaA => P(3)(63),lamdaB => P(3)(127),lamdaOut => P(2)(63));
G364: entity G port map(lamdaA => P(3)(0),lamdaB => P(3)(64),s => s(3)(0),lamdaOut => P(2)(64));
G365: entity G port map(lamdaA => P(3)(1),lamdaB => P(3)(65),s => s(3)(1),lamdaOut => P(2)(65));
G366: entity G port map(lamdaA => P(3)(2),lamdaB => P(3)(66),s => s(3)(2),lamdaOut => P(2)(66));
G367: entity G port map(lamdaA => P(3)(3),lamdaB => P(3)(67),s => s(3)(3),lamdaOut => P(2)(67));
G368: entity G port map(lamdaA => P(3)(4),lamdaB => P(3)(68),s => s(3)(4),lamdaOut => P(2)(68));
G369: entity G port map(lamdaA => P(3)(5),lamdaB => P(3)(69),s => s(3)(5),lamdaOut => P(2)(69));
G370: entity G port map(lamdaA => P(3)(6),lamdaB => P(3)(70),s => s(3)(6),lamdaOut => P(2)(70));
G371: entity G port map(lamdaA => P(3)(7),lamdaB => P(3)(71),s => s(3)(7),lamdaOut => P(2)(71));
G372: entity G port map(lamdaA => P(3)(8),lamdaB => P(3)(72),s => s(3)(8),lamdaOut => P(2)(72));
G373: entity G port map(lamdaA => P(3)(9),lamdaB => P(3)(73),s => s(3)(9),lamdaOut => P(2)(73));
G374: entity G port map(lamdaA => P(3)(10),lamdaB => P(3)(74),s => s(3)(10),lamdaOut => P(2)(74));
G375: entity G port map(lamdaA => P(3)(11),lamdaB => P(3)(75),s => s(3)(11),lamdaOut => P(2)(75));
G376: entity G port map(lamdaA => P(3)(12),lamdaB => P(3)(76),s => s(3)(12),lamdaOut => P(2)(76));
G377: entity G port map(lamdaA => P(3)(13),lamdaB => P(3)(77),s => s(3)(13),lamdaOut => P(2)(77));
G378: entity G port map(lamdaA => P(3)(14),lamdaB => P(3)(78),s => s(3)(14),lamdaOut => P(2)(78));
G379: entity G port map(lamdaA => P(3)(15),lamdaB => P(3)(79),s => s(3)(15),lamdaOut => P(2)(79));
G380: entity G port map(lamdaA => P(3)(16),lamdaB => P(3)(80),s => s(3)(16),lamdaOut => P(2)(80));
G381: entity G port map(lamdaA => P(3)(17),lamdaB => P(3)(81),s => s(3)(17),lamdaOut => P(2)(81));
G382: entity G port map(lamdaA => P(3)(18),lamdaB => P(3)(82),s => s(3)(18),lamdaOut => P(2)(82));
G383: entity G port map(lamdaA => P(3)(19),lamdaB => P(3)(83),s => s(3)(19),lamdaOut => P(2)(83));
G384: entity G port map(lamdaA => P(3)(20),lamdaB => P(3)(84),s => s(3)(20),lamdaOut => P(2)(84));
G385: entity G port map(lamdaA => P(3)(21),lamdaB => P(3)(85),s => s(3)(21),lamdaOut => P(2)(85));
G386: entity G port map(lamdaA => P(3)(22),lamdaB => P(3)(86),s => s(3)(22),lamdaOut => P(2)(86));
G387: entity G port map(lamdaA => P(3)(23),lamdaB => P(3)(87),s => s(3)(23),lamdaOut => P(2)(87));
G388: entity G port map(lamdaA => P(3)(24),lamdaB => P(3)(88),s => s(3)(24),lamdaOut => P(2)(88));
G389: entity G port map(lamdaA => P(3)(25),lamdaB => P(3)(89),s => s(3)(25),lamdaOut => P(2)(89));
G390: entity G port map(lamdaA => P(3)(26),lamdaB => P(3)(90),s => s(3)(26),lamdaOut => P(2)(90));
G391: entity G port map(lamdaA => P(3)(27),lamdaB => P(3)(91),s => s(3)(27),lamdaOut => P(2)(91));
G392: entity G port map(lamdaA => P(3)(28),lamdaB => P(3)(92),s => s(3)(28),lamdaOut => P(2)(92));
G393: entity G port map(lamdaA => P(3)(29),lamdaB => P(3)(93),s => s(3)(29),lamdaOut => P(2)(93));
G394: entity G port map(lamdaA => P(3)(30),lamdaB => P(3)(94),s => s(3)(30),lamdaOut => P(2)(94));
G395: entity G port map(lamdaA => P(3)(31),lamdaB => P(3)(95),s => s(3)(31),lamdaOut => P(2)(95));
G396: entity G port map(lamdaA => P(3)(32),lamdaB => P(3)(96),s => s(3)(32),lamdaOut => P(2)(96));
G397: entity G port map(lamdaA => P(3)(33),lamdaB => P(3)(97),s => s(3)(33),lamdaOut => P(2)(97));
G398: entity G port map(lamdaA => P(3)(34),lamdaB => P(3)(98),s => s(3)(34),lamdaOut => P(2)(98));
G399: entity G port map(lamdaA => P(3)(35),lamdaB => P(3)(99),s => s(3)(35),lamdaOut => P(2)(99));
G3100: entity G port map(lamdaA => P(3)(36),lamdaB => P(3)(100),s => s(3)(36),lamdaOut => P(2)(100));
G3101: entity G port map(lamdaA => P(3)(37),lamdaB => P(3)(101),s => s(3)(37),lamdaOut => P(2)(101));
G3102: entity G port map(lamdaA => P(3)(38),lamdaB => P(3)(102),s => s(3)(38),lamdaOut => P(2)(102));
G3103: entity G port map(lamdaA => P(3)(39),lamdaB => P(3)(103),s => s(3)(39),lamdaOut => P(2)(103));
G3104: entity G port map(lamdaA => P(3)(40),lamdaB => P(3)(104),s => s(3)(40),lamdaOut => P(2)(104));
G3105: entity G port map(lamdaA => P(3)(41),lamdaB => P(3)(105),s => s(3)(41),lamdaOut => P(2)(105));
G3106: entity G port map(lamdaA => P(3)(42),lamdaB => P(3)(106),s => s(3)(42),lamdaOut => P(2)(106));
G3107: entity G port map(lamdaA => P(3)(43),lamdaB => P(3)(107),s => s(3)(43),lamdaOut => P(2)(107));
G3108: entity G port map(lamdaA => P(3)(44),lamdaB => P(3)(108),s => s(3)(44),lamdaOut => P(2)(108));
G3109: entity G port map(lamdaA => P(3)(45),lamdaB => P(3)(109),s => s(3)(45),lamdaOut => P(2)(109));
G3110: entity G port map(lamdaA => P(3)(46),lamdaB => P(3)(110),s => s(3)(46),lamdaOut => P(2)(110));
G3111: entity G port map(lamdaA => P(3)(47),lamdaB => P(3)(111),s => s(3)(47),lamdaOut => P(2)(111));
G3112: entity G port map(lamdaA => P(3)(48),lamdaB => P(3)(112),s => s(3)(48),lamdaOut => P(2)(112));
G3113: entity G port map(lamdaA => P(3)(49),lamdaB => P(3)(113),s => s(3)(49),lamdaOut => P(2)(113));
G3114: entity G port map(lamdaA => P(3)(50),lamdaB => P(3)(114),s => s(3)(50),lamdaOut => P(2)(114));
G3115: entity G port map(lamdaA => P(3)(51),lamdaB => P(3)(115),s => s(3)(51),lamdaOut => P(2)(115));
G3116: entity G port map(lamdaA => P(3)(52),lamdaB => P(3)(116),s => s(3)(52),lamdaOut => P(2)(116));
G3117: entity G port map(lamdaA => P(3)(53),lamdaB => P(3)(117),s => s(3)(53),lamdaOut => P(2)(117));
G3118: entity G port map(lamdaA => P(3)(54),lamdaB => P(3)(118),s => s(3)(54),lamdaOut => P(2)(118));
G3119: entity G port map(lamdaA => P(3)(55),lamdaB => P(3)(119),s => s(3)(55),lamdaOut => P(2)(119));
G3120: entity G port map(lamdaA => P(3)(56),lamdaB => P(3)(120),s => s(3)(56),lamdaOut => P(2)(120));
G3121: entity G port map(lamdaA => P(3)(57),lamdaB => P(3)(121),s => s(3)(57),lamdaOut => P(2)(121));
G3122: entity G port map(lamdaA => P(3)(58),lamdaB => P(3)(122),s => s(3)(58),lamdaOut => P(2)(122));
G3123: entity G port map(lamdaA => P(3)(59),lamdaB => P(3)(123),s => s(3)(59),lamdaOut => P(2)(123));
G3124: entity G port map(lamdaA => P(3)(60),lamdaB => P(3)(124),s => s(3)(60),lamdaOut => P(2)(124));
G3125: entity G port map(lamdaA => P(3)(61),lamdaB => P(3)(125),s => s(3)(61),lamdaOut => P(2)(125));
G3126: entity G port map(lamdaA => P(3)(62),lamdaB => P(3)(126),s => s(3)(62),lamdaOut => P(2)(126));
G3127: entity G port map(lamdaA => P(3)(63),lamdaB => P(3)(127),s => s(3)(63),lamdaOut => P(2)(127));
F3128: entity F port map(lamdaA => P(3)(128),lamdaB => P(3)(192),lamdaOut => P(2)(128));
F3129: entity F port map(lamdaA => P(3)(129),lamdaB => P(3)(193),lamdaOut => P(2)(129));
F3130: entity F port map(lamdaA => P(3)(130),lamdaB => P(3)(194),lamdaOut => P(2)(130));
F3131: entity F port map(lamdaA => P(3)(131),lamdaB => P(3)(195),lamdaOut => P(2)(131));
F3132: entity F port map(lamdaA => P(3)(132),lamdaB => P(3)(196),lamdaOut => P(2)(132));
F3133: entity F port map(lamdaA => P(3)(133),lamdaB => P(3)(197),lamdaOut => P(2)(133));
F3134: entity F port map(lamdaA => P(3)(134),lamdaB => P(3)(198),lamdaOut => P(2)(134));
F3135: entity F port map(lamdaA => P(3)(135),lamdaB => P(3)(199),lamdaOut => P(2)(135));
F3136: entity F port map(lamdaA => P(3)(136),lamdaB => P(3)(200),lamdaOut => P(2)(136));
F3137: entity F port map(lamdaA => P(3)(137),lamdaB => P(3)(201),lamdaOut => P(2)(137));
F3138: entity F port map(lamdaA => P(3)(138),lamdaB => P(3)(202),lamdaOut => P(2)(138));
F3139: entity F port map(lamdaA => P(3)(139),lamdaB => P(3)(203),lamdaOut => P(2)(139));
F3140: entity F port map(lamdaA => P(3)(140),lamdaB => P(3)(204),lamdaOut => P(2)(140));
F3141: entity F port map(lamdaA => P(3)(141),lamdaB => P(3)(205),lamdaOut => P(2)(141));
F3142: entity F port map(lamdaA => P(3)(142),lamdaB => P(3)(206),lamdaOut => P(2)(142));
F3143: entity F port map(lamdaA => P(3)(143),lamdaB => P(3)(207),lamdaOut => P(2)(143));
F3144: entity F port map(lamdaA => P(3)(144),lamdaB => P(3)(208),lamdaOut => P(2)(144));
F3145: entity F port map(lamdaA => P(3)(145),lamdaB => P(3)(209),lamdaOut => P(2)(145));
F3146: entity F port map(lamdaA => P(3)(146),lamdaB => P(3)(210),lamdaOut => P(2)(146));
F3147: entity F port map(lamdaA => P(3)(147),lamdaB => P(3)(211),lamdaOut => P(2)(147));
F3148: entity F port map(lamdaA => P(3)(148),lamdaB => P(3)(212),lamdaOut => P(2)(148));
F3149: entity F port map(lamdaA => P(3)(149),lamdaB => P(3)(213),lamdaOut => P(2)(149));
F3150: entity F port map(lamdaA => P(3)(150),lamdaB => P(3)(214),lamdaOut => P(2)(150));
F3151: entity F port map(lamdaA => P(3)(151),lamdaB => P(3)(215),lamdaOut => P(2)(151));
F3152: entity F port map(lamdaA => P(3)(152),lamdaB => P(3)(216),lamdaOut => P(2)(152));
F3153: entity F port map(lamdaA => P(3)(153),lamdaB => P(3)(217),lamdaOut => P(2)(153));
F3154: entity F port map(lamdaA => P(3)(154),lamdaB => P(3)(218),lamdaOut => P(2)(154));
F3155: entity F port map(lamdaA => P(3)(155),lamdaB => P(3)(219),lamdaOut => P(2)(155));
F3156: entity F port map(lamdaA => P(3)(156),lamdaB => P(3)(220),lamdaOut => P(2)(156));
F3157: entity F port map(lamdaA => P(3)(157),lamdaB => P(3)(221),lamdaOut => P(2)(157));
F3158: entity F port map(lamdaA => P(3)(158),lamdaB => P(3)(222),lamdaOut => P(2)(158));
F3159: entity F port map(lamdaA => P(3)(159),lamdaB => P(3)(223),lamdaOut => P(2)(159));
F3160: entity F port map(lamdaA => P(3)(160),lamdaB => P(3)(224),lamdaOut => P(2)(160));
F3161: entity F port map(lamdaA => P(3)(161),lamdaB => P(3)(225),lamdaOut => P(2)(161));
F3162: entity F port map(lamdaA => P(3)(162),lamdaB => P(3)(226),lamdaOut => P(2)(162));
F3163: entity F port map(lamdaA => P(3)(163),lamdaB => P(3)(227),lamdaOut => P(2)(163));
F3164: entity F port map(lamdaA => P(3)(164),lamdaB => P(3)(228),lamdaOut => P(2)(164));
F3165: entity F port map(lamdaA => P(3)(165),lamdaB => P(3)(229),lamdaOut => P(2)(165));
F3166: entity F port map(lamdaA => P(3)(166),lamdaB => P(3)(230),lamdaOut => P(2)(166));
F3167: entity F port map(lamdaA => P(3)(167),lamdaB => P(3)(231),lamdaOut => P(2)(167));
F3168: entity F port map(lamdaA => P(3)(168),lamdaB => P(3)(232),lamdaOut => P(2)(168));
F3169: entity F port map(lamdaA => P(3)(169),lamdaB => P(3)(233),lamdaOut => P(2)(169));
F3170: entity F port map(lamdaA => P(3)(170),lamdaB => P(3)(234),lamdaOut => P(2)(170));
F3171: entity F port map(lamdaA => P(3)(171),lamdaB => P(3)(235),lamdaOut => P(2)(171));
F3172: entity F port map(lamdaA => P(3)(172),lamdaB => P(3)(236),lamdaOut => P(2)(172));
F3173: entity F port map(lamdaA => P(3)(173),lamdaB => P(3)(237),lamdaOut => P(2)(173));
F3174: entity F port map(lamdaA => P(3)(174),lamdaB => P(3)(238),lamdaOut => P(2)(174));
F3175: entity F port map(lamdaA => P(3)(175),lamdaB => P(3)(239),lamdaOut => P(2)(175));
F3176: entity F port map(lamdaA => P(3)(176),lamdaB => P(3)(240),lamdaOut => P(2)(176));
F3177: entity F port map(lamdaA => P(3)(177),lamdaB => P(3)(241),lamdaOut => P(2)(177));
F3178: entity F port map(lamdaA => P(3)(178),lamdaB => P(3)(242),lamdaOut => P(2)(178));
F3179: entity F port map(lamdaA => P(3)(179),lamdaB => P(3)(243),lamdaOut => P(2)(179));
F3180: entity F port map(lamdaA => P(3)(180),lamdaB => P(3)(244),lamdaOut => P(2)(180));
F3181: entity F port map(lamdaA => P(3)(181),lamdaB => P(3)(245),lamdaOut => P(2)(181));
F3182: entity F port map(lamdaA => P(3)(182),lamdaB => P(3)(246),lamdaOut => P(2)(182));
F3183: entity F port map(lamdaA => P(3)(183),lamdaB => P(3)(247),lamdaOut => P(2)(183));
F3184: entity F port map(lamdaA => P(3)(184),lamdaB => P(3)(248),lamdaOut => P(2)(184));
F3185: entity F port map(lamdaA => P(3)(185),lamdaB => P(3)(249),lamdaOut => P(2)(185));
F3186: entity F port map(lamdaA => P(3)(186),lamdaB => P(3)(250),lamdaOut => P(2)(186));
F3187: entity F port map(lamdaA => P(3)(187),lamdaB => P(3)(251),lamdaOut => P(2)(187));
F3188: entity F port map(lamdaA => P(3)(188),lamdaB => P(3)(252),lamdaOut => P(2)(188));
F3189: entity F port map(lamdaA => P(3)(189),lamdaB => P(3)(253),lamdaOut => P(2)(189));
F3190: entity F port map(lamdaA => P(3)(190),lamdaB => P(3)(254),lamdaOut => P(2)(190));
F3191: entity F port map(lamdaA => P(3)(191),lamdaB => P(3)(255),lamdaOut => P(2)(191));
G3192: entity G port map(lamdaA => P(3)(128),lamdaB => P(3)(192),s => s(3)(64),lamdaOut => P(2)(192));
G3193: entity G port map(lamdaA => P(3)(129),lamdaB => P(3)(193),s => s(3)(65),lamdaOut => P(2)(193));
G3194: entity G port map(lamdaA => P(3)(130),lamdaB => P(3)(194),s => s(3)(66),lamdaOut => P(2)(194));
G3195: entity G port map(lamdaA => P(3)(131),lamdaB => P(3)(195),s => s(3)(67),lamdaOut => P(2)(195));
G3196: entity G port map(lamdaA => P(3)(132),lamdaB => P(3)(196),s => s(3)(68),lamdaOut => P(2)(196));
G3197: entity G port map(lamdaA => P(3)(133),lamdaB => P(3)(197),s => s(3)(69),lamdaOut => P(2)(197));
G3198: entity G port map(lamdaA => P(3)(134),lamdaB => P(3)(198),s => s(3)(70),lamdaOut => P(2)(198));
G3199: entity G port map(lamdaA => P(3)(135),lamdaB => P(3)(199),s => s(3)(71),lamdaOut => P(2)(199));
G3200: entity G port map(lamdaA => P(3)(136),lamdaB => P(3)(200),s => s(3)(72),lamdaOut => P(2)(200));
G3201: entity G port map(lamdaA => P(3)(137),lamdaB => P(3)(201),s => s(3)(73),lamdaOut => P(2)(201));
G3202: entity G port map(lamdaA => P(3)(138),lamdaB => P(3)(202),s => s(3)(74),lamdaOut => P(2)(202));
G3203: entity G port map(lamdaA => P(3)(139),lamdaB => P(3)(203),s => s(3)(75),lamdaOut => P(2)(203));
G3204: entity G port map(lamdaA => P(3)(140),lamdaB => P(3)(204),s => s(3)(76),lamdaOut => P(2)(204));
G3205: entity G port map(lamdaA => P(3)(141),lamdaB => P(3)(205),s => s(3)(77),lamdaOut => P(2)(205));
G3206: entity G port map(lamdaA => P(3)(142),lamdaB => P(3)(206),s => s(3)(78),lamdaOut => P(2)(206));
G3207: entity G port map(lamdaA => P(3)(143),lamdaB => P(3)(207),s => s(3)(79),lamdaOut => P(2)(207));
G3208: entity G port map(lamdaA => P(3)(144),lamdaB => P(3)(208),s => s(3)(80),lamdaOut => P(2)(208));
G3209: entity G port map(lamdaA => P(3)(145),lamdaB => P(3)(209),s => s(3)(81),lamdaOut => P(2)(209));
G3210: entity G port map(lamdaA => P(3)(146),lamdaB => P(3)(210),s => s(3)(82),lamdaOut => P(2)(210));
G3211: entity G port map(lamdaA => P(3)(147),lamdaB => P(3)(211),s => s(3)(83),lamdaOut => P(2)(211));
G3212: entity G port map(lamdaA => P(3)(148),lamdaB => P(3)(212),s => s(3)(84),lamdaOut => P(2)(212));
G3213: entity G port map(lamdaA => P(3)(149),lamdaB => P(3)(213),s => s(3)(85),lamdaOut => P(2)(213));
G3214: entity G port map(lamdaA => P(3)(150),lamdaB => P(3)(214),s => s(3)(86),lamdaOut => P(2)(214));
G3215: entity G port map(lamdaA => P(3)(151),lamdaB => P(3)(215),s => s(3)(87),lamdaOut => P(2)(215));
G3216: entity G port map(lamdaA => P(3)(152),lamdaB => P(3)(216),s => s(3)(88),lamdaOut => P(2)(216));
G3217: entity G port map(lamdaA => P(3)(153),lamdaB => P(3)(217),s => s(3)(89),lamdaOut => P(2)(217));
G3218: entity G port map(lamdaA => P(3)(154),lamdaB => P(3)(218),s => s(3)(90),lamdaOut => P(2)(218));
G3219: entity G port map(lamdaA => P(3)(155),lamdaB => P(3)(219),s => s(3)(91),lamdaOut => P(2)(219));
G3220: entity G port map(lamdaA => P(3)(156),lamdaB => P(3)(220),s => s(3)(92),lamdaOut => P(2)(220));
G3221: entity G port map(lamdaA => P(3)(157),lamdaB => P(3)(221),s => s(3)(93),lamdaOut => P(2)(221));
G3222: entity G port map(lamdaA => P(3)(158),lamdaB => P(3)(222),s => s(3)(94),lamdaOut => P(2)(222));
G3223: entity G port map(lamdaA => P(3)(159),lamdaB => P(3)(223),s => s(3)(95),lamdaOut => P(2)(223));
G3224: entity G port map(lamdaA => P(3)(160),lamdaB => P(3)(224),s => s(3)(96),lamdaOut => P(2)(224));
G3225: entity G port map(lamdaA => P(3)(161),lamdaB => P(3)(225),s => s(3)(97),lamdaOut => P(2)(225));
G3226: entity G port map(lamdaA => P(3)(162),lamdaB => P(3)(226),s => s(3)(98),lamdaOut => P(2)(226));
G3227: entity G port map(lamdaA => P(3)(163),lamdaB => P(3)(227),s => s(3)(99),lamdaOut => P(2)(227));
G3228: entity G port map(lamdaA => P(3)(164),lamdaB => P(3)(228),s => s(3)(100),lamdaOut => P(2)(228));
G3229: entity G port map(lamdaA => P(3)(165),lamdaB => P(3)(229),s => s(3)(101),lamdaOut => P(2)(229));
G3230: entity G port map(lamdaA => P(3)(166),lamdaB => P(3)(230),s => s(3)(102),lamdaOut => P(2)(230));
G3231: entity G port map(lamdaA => P(3)(167),lamdaB => P(3)(231),s => s(3)(103),lamdaOut => P(2)(231));
G3232: entity G port map(lamdaA => P(3)(168),lamdaB => P(3)(232),s => s(3)(104),lamdaOut => P(2)(232));
G3233: entity G port map(lamdaA => P(3)(169),lamdaB => P(3)(233),s => s(3)(105),lamdaOut => P(2)(233));
G3234: entity G port map(lamdaA => P(3)(170),lamdaB => P(3)(234),s => s(3)(106),lamdaOut => P(2)(234));
G3235: entity G port map(lamdaA => P(3)(171),lamdaB => P(3)(235),s => s(3)(107),lamdaOut => P(2)(235));
G3236: entity G port map(lamdaA => P(3)(172),lamdaB => P(3)(236),s => s(3)(108),lamdaOut => P(2)(236));
G3237: entity G port map(lamdaA => P(3)(173),lamdaB => P(3)(237),s => s(3)(109),lamdaOut => P(2)(237));
G3238: entity G port map(lamdaA => P(3)(174),lamdaB => P(3)(238),s => s(3)(110),lamdaOut => P(2)(238));
G3239: entity G port map(lamdaA => P(3)(175),lamdaB => P(3)(239),s => s(3)(111),lamdaOut => P(2)(239));
G3240: entity G port map(lamdaA => P(3)(176),lamdaB => P(3)(240),s => s(3)(112),lamdaOut => P(2)(240));
G3241: entity G port map(lamdaA => P(3)(177),lamdaB => P(3)(241),s => s(3)(113),lamdaOut => P(2)(241));
G3242: entity G port map(lamdaA => P(3)(178),lamdaB => P(3)(242),s => s(3)(114),lamdaOut => P(2)(242));
G3243: entity G port map(lamdaA => P(3)(179),lamdaB => P(3)(243),s => s(3)(115),lamdaOut => P(2)(243));
G3244: entity G port map(lamdaA => P(3)(180),lamdaB => P(3)(244),s => s(3)(116),lamdaOut => P(2)(244));
G3245: entity G port map(lamdaA => P(3)(181),lamdaB => P(3)(245),s => s(3)(117),lamdaOut => P(2)(245));
G3246: entity G port map(lamdaA => P(3)(182),lamdaB => P(3)(246),s => s(3)(118),lamdaOut => P(2)(246));
G3247: entity G port map(lamdaA => P(3)(183),lamdaB => P(3)(247),s => s(3)(119),lamdaOut => P(2)(247));
G3248: entity G port map(lamdaA => P(3)(184),lamdaB => P(3)(248),s => s(3)(120),lamdaOut => P(2)(248));
G3249: entity G port map(lamdaA => P(3)(185),lamdaB => P(3)(249),s => s(3)(121),lamdaOut => P(2)(249));
G3250: entity G port map(lamdaA => P(3)(186),lamdaB => P(3)(250),s => s(3)(122),lamdaOut => P(2)(250));
G3251: entity G port map(lamdaA => P(3)(187),lamdaB => P(3)(251),s => s(3)(123),lamdaOut => P(2)(251));
G3252: entity G port map(lamdaA => P(3)(188),lamdaB => P(3)(252),s => s(3)(124),lamdaOut => P(2)(252));
G3253: entity G port map(lamdaA => P(3)(189),lamdaB => P(3)(253),s => s(3)(125),lamdaOut => P(2)(253));
G3254: entity G port map(lamdaA => P(3)(190),lamdaB => P(3)(254),s => s(3)(126),lamdaOut => P(2)(254));
G3255: entity G port map(lamdaA => P(3)(191),lamdaB => P(3)(255),s => s(3)(127),lamdaOut => P(2)(255));
F3256: entity F port map(lamdaA => P(3)(256),lamdaB => P(3)(320),lamdaOut => P(2)(256));
F3257: entity F port map(lamdaA => P(3)(257),lamdaB => P(3)(321),lamdaOut => P(2)(257));
F3258: entity F port map(lamdaA => P(3)(258),lamdaB => P(3)(322),lamdaOut => P(2)(258));
F3259: entity F port map(lamdaA => P(3)(259),lamdaB => P(3)(323),lamdaOut => P(2)(259));
F3260: entity F port map(lamdaA => P(3)(260),lamdaB => P(3)(324),lamdaOut => P(2)(260));
F3261: entity F port map(lamdaA => P(3)(261),lamdaB => P(3)(325),lamdaOut => P(2)(261));
F3262: entity F port map(lamdaA => P(3)(262),lamdaB => P(3)(326),lamdaOut => P(2)(262));
F3263: entity F port map(lamdaA => P(3)(263),lamdaB => P(3)(327),lamdaOut => P(2)(263));
F3264: entity F port map(lamdaA => P(3)(264),lamdaB => P(3)(328),lamdaOut => P(2)(264));
F3265: entity F port map(lamdaA => P(3)(265),lamdaB => P(3)(329),lamdaOut => P(2)(265));
F3266: entity F port map(lamdaA => P(3)(266),lamdaB => P(3)(330),lamdaOut => P(2)(266));
F3267: entity F port map(lamdaA => P(3)(267),lamdaB => P(3)(331),lamdaOut => P(2)(267));
F3268: entity F port map(lamdaA => P(3)(268),lamdaB => P(3)(332),lamdaOut => P(2)(268));
F3269: entity F port map(lamdaA => P(3)(269),lamdaB => P(3)(333),lamdaOut => P(2)(269));
F3270: entity F port map(lamdaA => P(3)(270),lamdaB => P(3)(334),lamdaOut => P(2)(270));
F3271: entity F port map(lamdaA => P(3)(271),lamdaB => P(3)(335),lamdaOut => P(2)(271));
F3272: entity F port map(lamdaA => P(3)(272),lamdaB => P(3)(336),lamdaOut => P(2)(272));
F3273: entity F port map(lamdaA => P(3)(273),lamdaB => P(3)(337),lamdaOut => P(2)(273));
F3274: entity F port map(lamdaA => P(3)(274),lamdaB => P(3)(338),lamdaOut => P(2)(274));
F3275: entity F port map(lamdaA => P(3)(275),lamdaB => P(3)(339),lamdaOut => P(2)(275));
F3276: entity F port map(lamdaA => P(3)(276),lamdaB => P(3)(340),lamdaOut => P(2)(276));
F3277: entity F port map(lamdaA => P(3)(277),lamdaB => P(3)(341),lamdaOut => P(2)(277));
F3278: entity F port map(lamdaA => P(3)(278),lamdaB => P(3)(342),lamdaOut => P(2)(278));
F3279: entity F port map(lamdaA => P(3)(279),lamdaB => P(3)(343),lamdaOut => P(2)(279));
F3280: entity F port map(lamdaA => P(3)(280),lamdaB => P(3)(344),lamdaOut => P(2)(280));
F3281: entity F port map(lamdaA => P(3)(281),lamdaB => P(3)(345),lamdaOut => P(2)(281));
F3282: entity F port map(lamdaA => P(3)(282),lamdaB => P(3)(346),lamdaOut => P(2)(282));
F3283: entity F port map(lamdaA => P(3)(283),lamdaB => P(3)(347),lamdaOut => P(2)(283));
F3284: entity F port map(lamdaA => P(3)(284),lamdaB => P(3)(348),lamdaOut => P(2)(284));
F3285: entity F port map(lamdaA => P(3)(285),lamdaB => P(3)(349),lamdaOut => P(2)(285));
F3286: entity F port map(lamdaA => P(3)(286),lamdaB => P(3)(350),lamdaOut => P(2)(286));
F3287: entity F port map(lamdaA => P(3)(287),lamdaB => P(3)(351),lamdaOut => P(2)(287));
F3288: entity F port map(lamdaA => P(3)(288),lamdaB => P(3)(352),lamdaOut => P(2)(288));
F3289: entity F port map(lamdaA => P(3)(289),lamdaB => P(3)(353),lamdaOut => P(2)(289));
F3290: entity F port map(lamdaA => P(3)(290),lamdaB => P(3)(354),lamdaOut => P(2)(290));
F3291: entity F port map(lamdaA => P(3)(291),lamdaB => P(3)(355),lamdaOut => P(2)(291));
F3292: entity F port map(lamdaA => P(3)(292),lamdaB => P(3)(356),lamdaOut => P(2)(292));
F3293: entity F port map(lamdaA => P(3)(293),lamdaB => P(3)(357),lamdaOut => P(2)(293));
F3294: entity F port map(lamdaA => P(3)(294),lamdaB => P(3)(358),lamdaOut => P(2)(294));
F3295: entity F port map(lamdaA => P(3)(295),lamdaB => P(3)(359),lamdaOut => P(2)(295));
F3296: entity F port map(lamdaA => P(3)(296),lamdaB => P(3)(360),lamdaOut => P(2)(296));
F3297: entity F port map(lamdaA => P(3)(297),lamdaB => P(3)(361),lamdaOut => P(2)(297));
F3298: entity F port map(lamdaA => P(3)(298),lamdaB => P(3)(362),lamdaOut => P(2)(298));
F3299: entity F port map(lamdaA => P(3)(299),lamdaB => P(3)(363),lamdaOut => P(2)(299));
F3300: entity F port map(lamdaA => P(3)(300),lamdaB => P(3)(364),lamdaOut => P(2)(300));
F3301: entity F port map(lamdaA => P(3)(301),lamdaB => P(3)(365),lamdaOut => P(2)(301));
F3302: entity F port map(lamdaA => P(3)(302),lamdaB => P(3)(366),lamdaOut => P(2)(302));
F3303: entity F port map(lamdaA => P(3)(303),lamdaB => P(3)(367),lamdaOut => P(2)(303));
F3304: entity F port map(lamdaA => P(3)(304),lamdaB => P(3)(368),lamdaOut => P(2)(304));
F3305: entity F port map(lamdaA => P(3)(305),lamdaB => P(3)(369),lamdaOut => P(2)(305));
F3306: entity F port map(lamdaA => P(3)(306),lamdaB => P(3)(370),lamdaOut => P(2)(306));
F3307: entity F port map(lamdaA => P(3)(307),lamdaB => P(3)(371),lamdaOut => P(2)(307));
F3308: entity F port map(lamdaA => P(3)(308),lamdaB => P(3)(372),lamdaOut => P(2)(308));
F3309: entity F port map(lamdaA => P(3)(309),lamdaB => P(3)(373),lamdaOut => P(2)(309));
F3310: entity F port map(lamdaA => P(3)(310),lamdaB => P(3)(374),lamdaOut => P(2)(310));
F3311: entity F port map(lamdaA => P(3)(311),lamdaB => P(3)(375),lamdaOut => P(2)(311));
F3312: entity F port map(lamdaA => P(3)(312),lamdaB => P(3)(376),lamdaOut => P(2)(312));
F3313: entity F port map(lamdaA => P(3)(313),lamdaB => P(3)(377),lamdaOut => P(2)(313));
F3314: entity F port map(lamdaA => P(3)(314),lamdaB => P(3)(378),lamdaOut => P(2)(314));
F3315: entity F port map(lamdaA => P(3)(315),lamdaB => P(3)(379),lamdaOut => P(2)(315));
F3316: entity F port map(lamdaA => P(3)(316),lamdaB => P(3)(380),lamdaOut => P(2)(316));
F3317: entity F port map(lamdaA => P(3)(317),lamdaB => P(3)(381),lamdaOut => P(2)(317));
F3318: entity F port map(lamdaA => P(3)(318),lamdaB => P(3)(382),lamdaOut => P(2)(318));
F3319: entity F port map(lamdaA => P(3)(319),lamdaB => P(3)(383),lamdaOut => P(2)(319));
G3320: entity G port map(lamdaA => P(3)(256),lamdaB => P(3)(320),s => s(3)(128),lamdaOut => P(2)(320));
G3321: entity G port map(lamdaA => P(3)(257),lamdaB => P(3)(321),s => s(3)(129),lamdaOut => P(2)(321));
G3322: entity G port map(lamdaA => P(3)(258),lamdaB => P(3)(322),s => s(3)(130),lamdaOut => P(2)(322));
G3323: entity G port map(lamdaA => P(3)(259),lamdaB => P(3)(323),s => s(3)(131),lamdaOut => P(2)(323));
G3324: entity G port map(lamdaA => P(3)(260),lamdaB => P(3)(324),s => s(3)(132),lamdaOut => P(2)(324));
G3325: entity G port map(lamdaA => P(3)(261),lamdaB => P(3)(325),s => s(3)(133),lamdaOut => P(2)(325));
G3326: entity G port map(lamdaA => P(3)(262),lamdaB => P(3)(326),s => s(3)(134),lamdaOut => P(2)(326));
G3327: entity G port map(lamdaA => P(3)(263),lamdaB => P(3)(327),s => s(3)(135),lamdaOut => P(2)(327));
G3328: entity G port map(lamdaA => P(3)(264),lamdaB => P(3)(328),s => s(3)(136),lamdaOut => P(2)(328));
G3329: entity G port map(lamdaA => P(3)(265),lamdaB => P(3)(329),s => s(3)(137),lamdaOut => P(2)(329));
G3330: entity G port map(lamdaA => P(3)(266),lamdaB => P(3)(330),s => s(3)(138),lamdaOut => P(2)(330));
G3331: entity G port map(lamdaA => P(3)(267),lamdaB => P(3)(331),s => s(3)(139),lamdaOut => P(2)(331));
G3332: entity G port map(lamdaA => P(3)(268),lamdaB => P(3)(332),s => s(3)(140),lamdaOut => P(2)(332));
G3333: entity G port map(lamdaA => P(3)(269),lamdaB => P(3)(333),s => s(3)(141),lamdaOut => P(2)(333));
G3334: entity G port map(lamdaA => P(3)(270),lamdaB => P(3)(334),s => s(3)(142),lamdaOut => P(2)(334));
G3335: entity G port map(lamdaA => P(3)(271),lamdaB => P(3)(335),s => s(3)(143),lamdaOut => P(2)(335));
G3336: entity G port map(lamdaA => P(3)(272),lamdaB => P(3)(336),s => s(3)(144),lamdaOut => P(2)(336));
G3337: entity G port map(lamdaA => P(3)(273),lamdaB => P(3)(337),s => s(3)(145),lamdaOut => P(2)(337));
G3338: entity G port map(lamdaA => P(3)(274),lamdaB => P(3)(338),s => s(3)(146),lamdaOut => P(2)(338));
G3339: entity G port map(lamdaA => P(3)(275),lamdaB => P(3)(339),s => s(3)(147),lamdaOut => P(2)(339));
G3340: entity G port map(lamdaA => P(3)(276),lamdaB => P(3)(340),s => s(3)(148),lamdaOut => P(2)(340));
G3341: entity G port map(lamdaA => P(3)(277),lamdaB => P(3)(341),s => s(3)(149),lamdaOut => P(2)(341));
G3342: entity G port map(lamdaA => P(3)(278),lamdaB => P(3)(342),s => s(3)(150),lamdaOut => P(2)(342));
G3343: entity G port map(lamdaA => P(3)(279),lamdaB => P(3)(343),s => s(3)(151),lamdaOut => P(2)(343));
G3344: entity G port map(lamdaA => P(3)(280),lamdaB => P(3)(344),s => s(3)(152),lamdaOut => P(2)(344));
G3345: entity G port map(lamdaA => P(3)(281),lamdaB => P(3)(345),s => s(3)(153),lamdaOut => P(2)(345));
G3346: entity G port map(lamdaA => P(3)(282),lamdaB => P(3)(346),s => s(3)(154),lamdaOut => P(2)(346));
G3347: entity G port map(lamdaA => P(3)(283),lamdaB => P(3)(347),s => s(3)(155),lamdaOut => P(2)(347));
G3348: entity G port map(lamdaA => P(3)(284),lamdaB => P(3)(348),s => s(3)(156),lamdaOut => P(2)(348));
G3349: entity G port map(lamdaA => P(3)(285),lamdaB => P(3)(349),s => s(3)(157),lamdaOut => P(2)(349));
G3350: entity G port map(lamdaA => P(3)(286),lamdaB => P(3)(350),s => s(3)(158),lamdaOut => P(2)(350));
G3351: entity G port map(lamdaA => P(3)(287),lamdaB => P(3)(351),s => s(3)(159),lamdaOut => P(2)(351));
G3352: entity G port map(lamdaA => P(3)(288),lamdaB => P(3)(352),s => s(3)(160),lamdaOut => P(2)(352));
G3353: entity G port map(lamdaA => P(3)(289),lamdaB => P(3)(353),s => s(3)(161),lamdaOut => P(2)(353));
G3354: entity G port map(lamdaA => P(3)(290),lamdaB => P(3)(354),s => s(3)(162),lamdaOut => P(2)(354));
G3355: entity G port map(lamdaA => P(3)(291),lamdaB => P(3)(355),s => s(3)(163),lamdaOut => P(2)(355));
G3356: entity G port map(lamdaA => P(3)(292),lamdaB => P(3)(356),s => s(3)(164),lamdaOut => P(2)(356));
G3357: entity G port map(lamdaA => P(3)(293),lamdaB => P(3)(357),s => s(3)(165),lamdaOut => P(2)(357));
G3358: entity G port map(lamdaA => P(3)(294),lamdaB => P(3)(358),s => s(3)(166),lamdaOut => P(2)(358));
G3359: entity G port map(lamdaA => P(3)(295),lamdaB => P(3)(359),s => s(3)(167),lamdaOut => P(2)(359));
G3360: entity G port map(lamdaA => P(3)(296),lamdaB => P(3)(360),s => s(3)(168),lamdaOut => P(2)(360));
G3361: entity G port map(lamdaA => P(3)(297),lamdaB => P(3)(361),s => s(3)(169),lamdaOut => P(2)(361));
G3362: entity G port map(lamdaA => P(3)(298),lamdaB => P(3)(362),s => s(3)(170),lamdaOut => P(2)(362));
G3363: entity G port map(lamdaA => P(3)(299),lamdaB => P(3)(363),s => s(3)(171),lamdaOut => P(2)(363));
G3364: entity G port map(lamdaA => P(3)(300),lamdaB => P(3)(364),s => s(3)(172),lamdaOut => P(2)(364));
G3365: entity G port map(lamdaA => P(3)(301),lamdaB => P(3)(365),s => s(3)(173),lamdaOut => P(2)(365));
G3366: entity G port map(lamdaA => P(3)(302),lamdaB => P(3)(366),s => s(3)(174),lamdaOut => P(2)(366));
G3367: entity G port map(lamdaA => P(3)(303),lamdaB => P(3)(367),s => s(3)(175),lamdaOut => P(2)(367));
G3368: entity G port map(lamdaA => P(3)(304),lamdaB => P(3)(368),s => s(3)(176),lamdaOut => P(2)(368));
G3369: entity G port map(lamdaA => P(3)(305),lamdaB => P(3)(369),s => s(3)(177),lamdaOut => P(2)(369));
G3370: entity G port map(lamdaA => P(3)(306),lamdaB => P(3)(370),s => s(3)(178),lamdaOut => P(2)(370));
G3371: entity G port map(lamdaA => P(3)(307),lamdaB => P(3)(371),s => s(3)(179),lamdaOut => P(2)(371));
G3372: entity G port map(lamdaA => P(3)(308),lamdaB => P(3)(372),s => s(3)(180),lamdaOut => P(2)(372));
G3373: entity G port map(lamdaA => P(3)(309),lamdaB => P(3)(373),s => s(3)(181),lamdaOut => P(2)(373));
G3374: entity G port map(lamdaA => P(3)(310),lamdaB => P(3)(374),s => s(3)(182),lamdaOut => P(2)(374));
G3375: entity G port map(lamdaA => P(3)(311),lamdaB => P(3)(375),s => s(3)(183),lamdaOut => P(2)(375));
G3376: entity G port map(lamdaA => P(3)(312),lamdaB => P(3)(376),s => s(3)(184),lamdaOut => P(2)(376));
G3377: entity G port map(lamdaA => P(3)(313),lamdaB => P(3)(377),s => s(3)(185),lamdaOut => P(2)(377));
G3378: entity G port map(lamdaA => P(3)(314),lamdaB => P(3)(378),s => s(3)(186),lamdaOut => P(2)(378));
G3379: entity G port map(lamdaA => P(3)(315),lamdaB => P(3)(379),s => s(3)(187),lamdaOut => P(2)(379));
G3380: entity G port map(lamdaA => P(3)(316),lamdaB => P(3)(380),s => s(3)(188),lamdaOut => P(2)(380));
G3381: entity G port map(lamdaA => P(3)(317),lamdaB => P(3)(381),s => s(3)(189),lamdaOut => P(2)(381));
G3382: entity G port map(lamdaA => P(3)(318),lamdaB => P(3)(382),s => s(3)(190),lamdaOut => P(2)(382));
G3383: entity G port map(lamdaA => P(3)(319),lamdaB => P(3)(383),s => s(3)(191),lamdaOut => P(2)(383));
F3384: entity F port map(lamdaA => P(3)(384),lamdaB => P(3)(448),lamdaOut => P(2)(384));
F3385: entity F port map(lamdaA => P(3)(385),lamdaB => P(3)(449),lamdaOut => P(2)(385));
F3386: entity F port map(lamdaA => P(3)(386),lamdaB => P(3)(450),lamdaOut => P(2)(386));
F3387: entity F port map(lamdaA => P(3)(387),lamdaB => P(3)(451),lamdaOut => P(2)(387));
F3388: entity F port map(lamdaA => P(3)(388),lamdaB => P(3)(452),lamdaOut => P(2)(388));
F3389: entity F port map(lamdaA => P(3)(389),lamdaB => P(3)(453),lamdaOut => P(2)(389));
F3390: entity F port map(lamdaA => P(3)(390),lamdaB => P(3)(454),lamdaOut => P(2)(390));
F3391: entity F port map(lamdaA => P(3)(391),lamdaB => P(3)(455),lamdaOut => P(2)(391));
F3392: entity F port map(lamdaA => P(3)(392),lamdaB => P(3)(456),lamdaOut => P(2)(392));
F3393: entity F port map(lamdaA => P(3)(393),lamdaB => P(3)(457),lamdaOut => P(2)(393));
F3394: entity F port map(lamdaA => P(3)(394),lamdaB => P(3)(458),lamdaOut => P(2)(394));
F3395: entity F port map(lamdaA => P(3)(395),lamdaB => P(3)(459),lamdaOut => P(2)(395));
F3396: entity F port map(lamdaA => P(3)(396),lamdaB => P(3)(460),lamdaOut => P(2)(396));
F3397: entity F port map(lamdaA => P(3)(397),lamdaB => P(3)(461),lamdaOut => P(2)(397));
F3398: entity F port map(lamdaA => P(3)(398),lamdaB => P(3)(462),lamdaOut => P(2)(398));
F3399: entity F port map(lamdaA => P(3)(399),lamdaB => P(3)(463),lamdaOut => P(2)(399));
F3400: entity F port map(lamdaA => P(3)(400),lamdaB => P(3)(464),lamdaOut => P(2)(400));
F3401: entity F port map(lamdaA => P(3)(401),lamdaB => P(3)(465),lamdaOut => P(2)(401));
F3402: entity F port map(lamdaA => P(3)(402),lamdaB => P(3)(466),lamdaOut => P(2)(402));
F3403: entity F port map(lamdaA => P(3)(403),lamdaB => P(3)(467),lamdaOut => P(2)(403));
F3404: entity F port map(lamdaA => P(3)(404),lamdaB => P(3)(468),lamdaOut => P(2)(404));
F3405: entity F port map(lamdaA => P(3)(405),lamdaB => P(3)(469),lamdaOut => P(2)(405));
F3406: entity F port map(lamdaA => P(3)(406),lamdaB => P(3)(470),lamdaOut => P(2)(406));
F3407: entity F port map(lamdaA => P(3)(407),lamdaB => P(3)(471),lamdaOut => P(2)(407));
F3408: entity F port map(lamdaA => P(3)(408),lamdaB => P(3)(472),lamdaOut => P(2)(408));
F3409: entity F port map(lamdaA => P(3)(409),lamdaB => P(3)(473),lamdaOut => P(2)(409));
F3410: entity F port map(lamdaA => P(3)(410),lamdaB => P(3)(474),lamdaOut => P(2)(410));
F3411: entity F port map(lamdaA => P(3)(411),lamdaB => P(3)(475),lamdaOut => P(2)(411));
F3412: entity F port map(lamdaA => P(3)(412),lamdaB => P(3)(476),lamdaOut => P(2)(412));
F3413: entity F port map(lamdaA => P(3)(413),lamdaB => P(3)(477),lamdaOut => P(2)(413));
F3414: entity F port map(lamdaA => P(3)(414),lamdaB => P(3)(478),lamdaOut => P(2)(414));
F3415: entity F port map(lamdaA => P(3)(415),lamdaB => P(3)(479),lamdaOut => P(2)(415));
F3416: entity F port map(lamdaA => P(3)(416),lamdaB => P(3)(480),lamdaOut => P(2)(416));
F3417: entity F port map(lamdaA => P(3)(417),lamdaB => P(3)(481),lamdaOut => P(2)(417));
F3418: entity F port map(lamdaA => P(3)(418),lamdaB => P(3)(482),lamdaOut => P(2)(418));
F3419: entity F port map(lamdaA => P(3)(419),lamdaB => P(3)(483),lamdaOut => P(2)(419));
F3420: entity F port map(lamdaA => P(3)(420),lamdaB => P(3)(484),lamdaOut => P(2)(420));
F3421: entity F port map(lamdaA => P(3)(421),lamdaB => P(3)(485),lamdaOut => P(2)(421));
F3422: entity F port map(lamdaA => P(3)(422),lamdaB => P(3)(486),lamdaOut => P(2)(422));
F3423: entity F port map(lamdaA => P(3)(423),lamdaB => P(3)(487),lamdaOut => P(2)(423));
F3424: entity F port map(lamdaA => P(3)(424),lamdaB => P(3)(488),lamdaOut => P(2)(424));
F3425: entity F port map(lamdaA => P(3)(425),lamdaB => P(3)(489),lamdaOut => P(2)(425));
F3426: entity F port map(lamdaA => P(3)(426),lamdaB => P(3)(490),lamdaOut => P(2)(426));
F3427: entity F port map(lamdaA => P(3)(427),lamdaB => P(3)(491),lamdaOut => P(2)(427));
F3428: entity F port map(lamdaA => P(3)(428),lamdaB => P(3)(492),lamdaOut => P(2)(428));
F3429: entity F port map(lamdaA => P(3)(429),lamdaB => P(3)(493),lamdaOut => P(2)(429));
F3430: entity F port map(lamdaA => P(3)(430),lamdaB => P(3)(494),lamdaOut => P(2)(430));
F3431: entity F port map(lamdaA => P(3)(431),lamdaB => P(3)(495),lamdaOut => P(2)(431));
F3432: entity F port map(lamdaA => P(3)(432),lamdaB => P(3)(496),lamdaOut => P(2)(432));
F3433: entity F port map(lamdaA => P(3)(433),lamdaB => P(3)(497),lamdaOut => P(2)(433));
F3434: entity F port map(lamdaA => P(3)(434),lamdaB => P(3)(498),lamdaOut => P(2)(434));
F3435: entity F port map(lamdaA => P(3)(435),lamdaB => P(3)(499),lamdaOut => P(2)(435));
F3436: entity F port map(lamdaA => P(3)(436),lamdaB => P(3)(500),lamdaOut => P(2)(436));
F3437: entity F port map(lamdaA => P(3)(437),lamdaB => P(3)(501),lamdaOut => P(2)(437));
F3438: entity F port map(lamdaA => P(3)(438),lamdaB => P(3)(502),lamdaOut => P(2)(438));
F3439: entity F port map(lamdaA => P(3)(439),lamdaB => P(3)(503),lamdaOut => P(2)(439));
F3440: entity F port map(lamdaA => P(3)(440),lamdaB => P(3)(504),lamdaOut => P(2)(440));
F3441: entity F port map(lamdaA => P(3)(441),lamdaB => P(3)(505),lamdaOut => P(2)(441));
F3442: entity F port map(lamdaA => P(3)(442),lamdaB => P(3)(506),lamdaOut => P(2)(442));
F3443: entity F port map(lamdaA => P(3)(443),lamdaB => P(3)(507),lamdaOut => P(2)(443));
F3444: entity F port map(lamdaA => P(3)(444),lamdaB => P(3)(508),lamdaOut => P(2)(444));
F3445: entity F port map(lamdaA => P(3)(445),lamdaB => P(3)(509),lamdaOut => P(2)(445));
F3446: entity F port map(lamdaA => P(3)(446),lamdaB => P(3)(510),lamdaOut => P(2)(446));
F3447: entity F port map(lamdaA => P(3)(447),lamdaB => P(3)(511),lamdaOut => P(2)(447));
G3448: entity G port map(lamdaA => P(3)(384),lamdaB => P(3)(448),s => s(3)(192),lamdaOut => P(2)(448));
G3449: entity G port map(lamdaA => P(3)(385),lamdaB => P(3)(449),s => s(3)(193),lamdaOut => P(2)(449));
G3450: entity G port map(lamdaA => P(3)(386),lamdaB => P(3)(450),s => s(3)(194),lamdaOut => P(2)(450));
G3451: entity G port map(lamdaA => P(3)(387),lamdaB => P(3)(451),s => s(3)(195),lamdaOut => P(2)(451));
G3452: entity G port map(lamdaA => P(3)(388),lamdaB => P(3)(452),s => s(3)(196),lamdaOut => P(2)(452));
G3453: entity G port map(lamdaA => P(3)(389),lamdaB => P(3)(453),s => s(3)(197),lamdaOut => P(2)(453));
G3454: entity G port map(lamdaA => P(3)(390),lamdaB => P(3)(454),s => s(3)(198),lamdaOut => P(2)(454));
G3455: entity G port map(lamdaA => P(3)(391),lamdaB => P(3)(455),s => s(3)(199),lamdaOut => P(2)(455));
G3456: entity G port map(lamdaA => P(3)(392),lamdaB => P(3)(456),s => s(3)(200),lamdaOut => P(2)(456));
G3457: entity G port map(lamdaA => P(3)(393),lamdaB => P(3)(457),s => s(3)(201),lamdaOut => P(2)(457));
G3458: entity G port map(lamdaA => P(3)(394),lamdaB => P(3)(458),s => s(3)(202),lamdaOut => P(2)(458));
G3459: entity G port map(lamdaA => P(3)(395),lamdaB => P(3)(459),s => s(3)(203),lamdaOut => P(2)(459));
G3460: entity G port map(lamdaA => P(3)(396),lamdaB => P(3)(460),s => s(3)(204),lamdaOut => P(2)(460));
G3461: entity G port map(lamdaA => P(3)(397),lamdaB => P(3)(461),s => s(3)(205),lamdaOut => P(2)(461));
G3462: entity G port map(lamdaA => P(3)(398),lamdaB => P(3)(462),s => s(3)(206),lamdaOut => P(2)(462));
G3463: entity G port map(lamdaA => P(3)(399),lamdaB => P(3)(463),s => s(3)(207),lamdaOut => P(2)(463));
G3464: entity G port map(lamdaA => P(3)(400),lamdaB => P(3)(464),s => s(3)(208),lamdaOut => P(2)(464));
G3465: entity G port map(lamdaA => P(3)(401),lamdaB => P(3)(465),s => s(3)(209),lamdaOut => P(2)(465));
G3466: entity G port map(lamdaA => P(3)(402),lamdaB => P(3)(466),s => s(3)(210),lamdaOut => P(2)(466));
G3467: entity G port map(lamdaA => P(3)(403),lamdaB => P(3)(467),s => s(3)(211),lamdaOut => P(2)(467));
G3468: entity G port map(lamdaA => P(3)(404),lamdaB => P(3)(468),s => s(3)(212),lamdaOut => P(2)(468));
G3469: entity G port map(lamdaA => P(3)(405),lamdaB => P(3)(469),s => s(3)(213),lamdaOut => P(2)(469));
G3470: entity G port map(lamdaA => P(3)(406),lamdaB => P(3)(470),s => s(3)(214),lamdaOut => P(2)(470));
G3471: entity G port map(lamdaA => P(3)(407),lamdaB => P(3)(471),s => s(3)(215),lamdaOut => P(2)(471));
G3472: entity G port map(lamdaA => P(3)(408),lamdaB => P(3)(472),s => s(3)(216),lamdaOut => P(2)(472));
G3473: entity G port map(lamdaA => P(3)(409),lamdaB => P(3)(473),s => s(3)(217),lamdaOut => P(2)(473));
G3474: entity G port map(lamdaA => P(3)(410),lamdaB => P(3)(474),s => s(3)(218),lamdaOut => P(2)(474));
G3475: entity G port map(lamdaA => P(3)(411),lamdaB => P(3)(475),s => s(3)(219),lamdaOut => P(2)(475));
G3476: entity G port map(lamdaA => P(3)(412),lamdaB => P(3)(476),s => s(3)(220),lamdaOut => P(2)(476));
G3477: entity G port map(lamdaA => P(3)(413),lamdaB => P(3)(477),s => s(3)(221),lamdaOut => P(2)(477));
G3478: entity G port map(lamdaA => P(3)(414),lamdaB => P(3)(478),s => s(3)(222),lamdaOut => P(2)(478));
G3479: entity G port map(lamdaA => P(3)(415),lamdaB => P(3)(479),s => s(3)(223),lamdaOut => P(2)(479));
G3480: entity G port map(lamdaA => P(3)(416),lamdaB => P(3)(480),s => s(3)(224),lamdaOut => P(2)(480));
G3481: entity G port map(lamdaA => P(3)(417),lamdaB => P(3)(481),s => s(3)(225),lamdaOut => P(2)(481));
G3482: entity G port map(lamdaA => P(3)(418),lamdaB => P(3)(482),s => s(3)(226),lamdaOut => P(2)(482));
G3483: entity G port map(lamdaA => P(3)(419),lamdaB => P(3)(483),s => s(3)(227),lamdaOut => P(2)(483));
G3484: entity G port map(lamdaA => P(3)(420),lamdaB => P(3)(484),s => s(3)(228),lamdaOut => P(2)(484));
G3485: entity G port map(lamdaA => P(3)(421),lamdaB => P(3)(485),s => s(3)(229),lamdaOut => P(2)(485));
G3486: entity G port map(lamdaA => P(3)(422),lamdaB => P(3)(486),s => s(3)(230),lamdaOut => P(2)(486));
G3487: entity G port map(lamdaA => P(3)(423),lamdaB => P(3)(487),s => s(3)(231),lamdaOut => P(2)(487));
G3488: entity G port map(lamdaA => P(3)(424),lamdaB => P(3)(488),s => s(3)(232),lamdaOut => P(2)(488));
G3489: entity G port map(lamdaA => P(3)(425),lamdaB => P(3)(489),s => s(3)(233),lamdaOut => P(2)(489));
G3490: entity G port map(lamdaA => P(3)(426),lamdaB => P(3)(490),s => s(3)(234),lamdaOut => P(2)(490));
G3491: entity G port map(lamdaA => P(3)(427),lamdaB => P(3)(491),s => s(3)(235),lamdaOut => P(2)(491));
G3492: entity G port map(lamdaA => P(3)(428),lamdaB => P(3)(492),s => s(3)(236),lamdaOut => P(2)(492));
G3493: entity G port map(lamdaA => P(3)(429),lamdaB => P(3)(493),s => s(3)(237),lamdaOut => P(2)(493));
G3494: entity G port map(lamdaA => P(3)(430),lamdaB => P(3)(494),s => s(3)(238),lamdaOut => P(2)(494));
G3495: entity G port map(lamdaA => P(3)(431),lamdaB => P(3)(495),s => s(3)(239),lamdaOut => P(2)(495));
G3496: entity G port map(lamdaA => P(3)(432),lamdaB => P(3)(496),s => s(3)(240),lamdaOut => P(2)(496));
G3497: entity G port map(lamdaA => P(3)(433),lamdaB => P(3)(497),s => s(3)(241),lamdaOut => P(2)(497));
G3498: entity G port map(lamdaA => P(3)(434),lamdaB => P(3)(498),s => s(3)(242),lamdaOut => P(2)(498));
G3499: entity G port map(lamdaA => P(3)(435),lamdaB => P(3)(499),s => s(3)(243),lamdaOut => P(2)(499));
G3500: entity G port map(lamdaA => P(3)(436),lamdaB => P(3)(500),s => s(3)(244),lamdaOut => P(2)(500));
G3501: entity G port map(lamdaA => P(3)(437),lamdaB => P(3)(501),s => s(3)(245),lamdaOut => P(2)(501));
G3502: entity G port map(lamdaA => P(3)(438),lamdaB => P(3)(502),s => s(3)(246),lamdaOut => P(2)(502));
G3503: entity G port map(lamdaA => P(3)(439),lamdaB => P(3)(503),s => s(3)(247),lamdaOut => P(2)(503));
G3504: entity G port map(lamdaA => P(3)(440),lamdaB => P(3)(504),s => s(3)(248),lamdaOut => P(2)(504));
G3505: entity G port map(lamdaA => P(3)(441),lamdaB => P(3)(505),s => s(3)(249),lamdaOut => P(2)(505));
G3506: entity G port map(lamdaA => P(3)(442),lamdaB => P(3)(506),s => s(3)(250),lamdaOut => P(2)(506));
G3507: entity G port map(lamdaA => P(3)(443),lamdaB => P(3)(507),s => s(3)(251),lamdaOut => P(2)(507));
G3508: entity G port map(lamdaA => P(3)(444),lamdaB => P(3)(508),s => s(3)(252),lamdaOut => P(2)(508));
G3509: entity G port map(lamdaA => P(3)(445),lamdaB => P(3)(509),s => s(3)(253),lamdaOut => P(2)(509));
G3510: entity G port map(lamdaA => P(3)(446),lamdaB => P(3)(510),s => s(3)(254),lamdaOut => P(2)(510));
G3511: entity G port map(lamdaA => P(3)(447),lamdaB => P(3)(511),s => s(3)(255),lamdaOut => P(2)(511));
-- STAGE 2
F20: entity F port map(lamdaA => P(2)(0),lamdaB => P(2)(128),lamdaOut => P(1)(0));
F21: entity F port map(lamdaA => P(2)(1),lamdaB => P(2)(129),lamdaOut => P(1)(1));
F22: entity F port map(lamdaA => P(2)(2),lamdaB => P(2)(130),lamdaOut => P(1)(2));
F23: entity F port map(lamdaA => P(2)(3),lamdaB => P(2)(131),lamdaOut => P(1)(3));
F24: entity F port map(lamdaA => P(2)(4),lamdaB => P(2)(132),lamdaOut => P(1)(4));
F25: entity F port map(lamdaA => P(2)(5),lamdaB => P(2)(133),lamdaOut => P(1)(5));
F26: entity F port map(lamdaA => P(2)(6),lamdaB => P(2)(134),lamdaOut => P(1)(6));
F27: entity F port map(lamdaA => P(2)(7),lamdaB => P(2)(135),lamdaOut => P(1)(7));
F28: entity F port map(lamdaA => P(2)(8),lamdaB => P(2)(136),lamdaOut => P(1)(8));
F29: entity F port map(lamdaA => P(2)(9),lamdaB => P(2)(137),lamdaOut => P(1)(9));
F210: entity F port map(lamdaA => P(2)(10),lamdaB => P(2)(138),lamdaOut => P(1)(10));
F211: entity F port map(lamdaA => P(2)(11),lamdaB => P(2)(139),lamdaOut => P(1)(11));
F212: entity F port map(lamdaA => P(2)(12),lamdaB => P(2)(140),lamdaOut => P(1)(12));
F213: entity F port map(lamdaA => P(2)(13),lamdaB => P(2)(141),lamdaOut => P(1)(13));
F214: entity F port map(lamdaA => P(2)(14),lamdaB => P(2)(142),lamdaOut => P(1)(14));
F215: entity F port map(lamdaA => P(2)(15),lamdaB => P(2)(143),lamdaOut => P(1)(15));
F216: entity F port map(lamdaA => P(2)(16),lamdaB => P(2)(144),lamdaOut => P(1)(16));
F217: entity F port map(lamdaA => P(2)(17),lamdaB => P(2)(145),lamdaOut => P(1)(17));
F218: entity F port map(lamdaA => P(2)(18),lamdaB => P(2)(146),lamdaOut => P(1)(18));
F219: entity F port map(lamdaA => P(2)(19),lamdaB => P(2)(147),lamdaOut => P(1)(19));
F220: entity F port map(lamdaA => P(2)(20),lamdaB => P(2)(148),lamdaOut => P(1)(20));
F221: entity F port map(lamdaA => P(2)(21),lamdaB => P(2)(149),lamdaOut => P(1)(21));
F222: entity F port map(lamdaA => P(2)(22),lamdaB => P(2)(150),lamdaOut => P(1)(22));
F223: entity F port map(lamdaA => P(2)(23),lamdaB => P(2)(151),lamdaOut => P(1)(23));
F224: entity F port map(lamdaA => P(2)(24),lamdaB => P(2)(152),lamdaOut => P(1)(24));
F225: entity F port map(lamdaA => P(2)(25),lamdaB => P(2)(153),lamdaOut => P(1)(25));
F226: entity F port map(lamdaA => P(2)(26),lamdaB => P(2)(154),lamdaOut => P(1)(26));
F227: entity F port map(lamdaA => P(2)(27),lamdaB => P(2)(155),lamdaOut => P(1)(27));
F228: entity F port map(lamdaA => P(2)(28),lamdaB => P(2)(156),lamdaOut => P(1)(28));
F229: entity F port map(lamdaA => P(2)(29),lamdaB => P(2)(157),lamdaOut => P(1)(29));
F230: entity F port map(lamdaA => P(2)(30),lamdaB => P(2)(158),lamdaOut => P(1)(30));
F231: entity F port map(lamdaA => P(2)(31),lamdaB => P(2)(159),lamdaOut => P(1)(31));
F232: entity F port map(lamdaA => P(2)(32),lamdaB => P(2)(160),lamdaOut => P(1)(32));
F233: entity F port map(lamdaA => P(2)(33),lamdaB => P(2)(161),lamdaOut => P(1)(33));
F234: entity F port map(lamdaA => P(2)(34),lamdaB => P(2)(162),lamdaOut => P(1)(34));
F235: entity F port map(lamdaA => P(2)(35),lamdaB => P(2)(163),lamdaOut => P(1)(35));
F236: entity F port map(lamdaA => P(2)(36),lamdaB => P(2)(164),lamdaOut => P(1)(36));
F237: entity F port map(lamdaA => P(2)(37),lamdaB => P(2)(165),lamdaOut => P(1)(37));
F238: entity F port map(lamdaA => P(2)(38),lamdaB => P(2)(166),lamdaOut => P(1)(38));
F239: entity F port map(lamdaA => P(2)(39),lamdaB => P(2)(167),lamdaOut => P(1)(39));
F240: entity F port map(lamdaA => P(2)(40),lamdaB => P(2)(168),lamdaOut => P(1)(40));
F241: entity F port map(lamdaA => P(2)(41),lamdaB => P(2)(169),lamdaOut => P(1)(41));
F242: entity F port map(lamdaA => P(2)(42),lamdaB => P(2)(170),lamdaOut => P(1)(42));
F243: entity F port map(lamdaA => P(2)(43),lamdaB => P(2)(171),lamdaOut => P(1)(43));
F244: entity F port map(lamdaA => P(2)(44),lamdaB => P(2)(172),lamdaOut => P(1)(44));
F245: entity F port map(lamdaA => P(2)(45),lamdaB => P(2)(173),lamdaOut => P(1)(45));
F246: entity F port map(lamdaA => P(2)(46),lamdaB => P(2)(174),lamdaOut => P(1)(46));
F247: entity F port map(lamdaA => P(2)(47),lamdaB => P(2)(175),lamdaOut => P(1)(47));
F248: entity F port map(lamdaA => P(2)(48),lamdaB => P(2)(176),lamdaOut => P(1)(48));
F249: entity F port map(lamdaA => P(2)(49),lamdaB => P(2)(177),lamdaOut => P(1)(49));
F250: entity F port map(lamdaA => P(2)(50),lamdaB => P(2)(178),lamdaOut => P(1)(50));
F251: entity F port map(lamdaA => P(2)(51),lamdaB => P(2)(179),lamdaOut => P(1)(51));
F252: entity F port map(lamdaA => P(2)(52),lamdaB => P(2)(180),lamdaOut => P(1)(52));
F253: entity F port map(lamdaA => P(2)(53),lamdaB => P(2)(181),lamdaOut => P(1)(53));
F254: entity F port map(lamdaA => P(2)(54),lamdaB => P(2)(182),lamdaOut => P(1)(54));
F255: entity F port map(lamdaA => P(2)(55),lamdaB => P(2)(183),lamdaOut => P(1)(55));
F256: entity F port map(lamdaA => P(2)(56),lamdaB => P(2)(184),lamdaOut => P(1)(56));
F257: entity F port map(lamdaA => P(2)(57),lamdaB => P(2)(185),lamdaOut => P(1)(57));
F258: entity F port map(lamdaA => P(2)(58),lamdaB => P(2)(186),lamdaOut => P(1)(58));
F259: entity F port map(lamdaA => P(2)(59),lamdaB => P(2)(187),lamdaOut => P(1)(59));
F260: entity F port map(lamdaA => P(2)(60),lamdaB => P(2)(188),lamdaOut => P(1)(60));
F261: entity F port map(lamdaA => P(2)(61),lamdaB => P(2)(189),lamdaOut => P(1)(61));
F262: entity F port map(lamdaA => P(2)(62),lamdaB => P(2)(190),lamdaOut => P(1)(62));
F263: entity F port map(lamdaA => P(2)(63),lamdaB => P(2)(191),lamdaOut => P(1)(63));
F264: entity F port map(lamdaA => P(2)(64),lamdaB => P(2)(192),lamdaOut => P(1)(64));
F265: entity F port map(lamdaA => P(2)(65),lamdaB => P(2)(193),lamdaOut => P(1)(65));
F266: entity F port map(lamdaA => P(2)(66),lamdaB => P(2)(194),lamdaOut => P(1)(66));
F267: entity F port map(lamdaA => P(2)(67),lamdaB => P(2)(195),lamdaOut => P(1)(67));
F268: entity F port map(lamdaA => P(2)(68),lamdaB => P(2)(196),lamdaOut => P(1)(68));
F269: entity F port map(lamdaA => P(2)(69),lamdaB => P(2)(197),lamdaOut => P(1)(69));
F270: entity F port map(lamdaA => P(2)(70),lamdaB => P(2)(198),lamdaOut => P(1)(70));
F271: entity F port map(lamdaA => P(2)(71),lamdaB => P(2)(199),lamdaOut => P(1)(71));
F272: entity F port map(lamdaA => P(2)(72),lamdaB => P(2)(200),lamdaOut => P(1)(72));
F273: entity F port map(lamdaA => P(2)(73),lamdaB => P(2)(201),lamdaOut => P(1)(73));
F274: entity F port map(lamdaA => P(2)(74),lamdaB => P(2)(202),lamdaOut => P(1)(74));
F275: entity F port map(lamdaA => P(2)(75),lamdaB => P(2)(203),lamdaOut => P(1)(75));
F276: entity F port map(lamdaA => P(2)(76),lamdaB => P(2)(204),lamdaOut => P(1)(76));
F277: entity F port map(lamdaA => P(2)(77),lamdaB => P(2)(205),lamdaOut => P(1)(77));
F278: entity F port map(lamdaA => P(2)(78),lamdaB => P(2)(206),lamdaOut => P(1)(78));
F279: entity F port map(lamdaA => P(2)(79),lamdaB => P(2)(207),lamdaOut => P(1)(79));
F280: entity F port map(lamdaA => P(2)(80),lamdaB => P(2)(208),lamdaOut => P(1)(80));
F281: entity F port map(lamdaA => P(2)(81),lamdaB => P(2)(209),lamdaOut => P(1)(81));
F282: entity F port map(lamdaA => P(2)(82),lamdaB => P(2)(210),lamdaOut => P(1)(82));
F283: entity F port map(lamdaA => P(2)(83),lamdaB => P(2)(211),lamdaOut => P(1)(83));
F284: entity F port map(lamdaA => P(2)(84),lamdaB => P(2)(212),lamdaOut => P(1)(84));
F285: entity F port map(lamdaA => P(2)(85),lamdaB => P(2)(213),lamdaOut => P(1)(85));
F286: entity F port map(lamdaA => P(2)(86),lamdaB => P(2)(214),lamdaOut => P(1)(86));
F287: entity F port map(lamdaA => P(2)(87),lamdaB => P(2)(215),lamdaOut => P(1)(87));
F288: entity F port map(lamdaA => P(2)(88),lamdaB => P(2)(216),lamdaOut => P(1)(88));
F289: entity F port map(lamdaA => P(2)(89),lamdaB => P(2)(217),lamdaOut => P(1)(89));
F290: entity F port map(lamdaA => P(2)(90),lamdaB => P(2)(218),lamdaOut => P(1)(90));
F291: entity F port map(lamdaA => P(2)(91),lamdaB => P(2)(219),lamdaOut => P(1)(91));
F292: entity F port map(lamdaA => P(2)(92),lamdaB => P(2)(220),lamdaOut => P(1)(92));
F293: entity F port map(lamdaA => P(2)(93),lamdaB => P(2)(221),lamdaOut => P(1)(93));
F294: entity F port map(lamdaA => P(2)(94),lamdaB => P(2)(222),lamdaOut => P(1)(94));
F295: entity F port map(lamdaA => P(2)(95),lamdaB => P(2)(223),lamdaOut => P(1)(95));
F296: entity F port map(lamdaA => P(2)(96),lamdaB => P(2)(224),lamdaOut => P(1)(96));
F297: entity F port map(lamdaA => P(2)(97),lamdaB => P(2)(225),lamdaOut => P(1)(97));
F298: entity F port map(lamdaA => P(2)(98),lamdaB => P(2)(226),lamdaOut => P(1)(98));
F299: entity F port map(lamdaA => P(2)(99),lamdaB => P(2)(227),lamdaOut => P(1)(99));
F2100: entity F port map(lamdaA => P(2)(100),lamdaB => P(2)(228),lamdaOut => P(1)(100));
F2101: entity F port map(lamdaA => P(2)(101),lamdaB => P(2)(229),lamdaOut => P(1)(101));
F2102: entity F port map(lamdaA => P(2)(102),lamdaB => P(2)(230),lamdaOut => P(1)(102));
F2103: entity F port map(lamdaA => P(2)(103),lamdaB => P(2)(231),lamdaOut => P(1)(103));
F2104: entity F port map(lamdaA => P(2)(104),lamdaB => P(2)(232),lamdaOut => P(1)(104));
F2105: entity F port map(lamdaA => P(2)(105),lamdaB => P(2)(233),lamdaOut => P(1)(105));
F2106: entity F port map(lamdaA => P(2)(106),lamdaB => P(2)(234),lamdaOut => P(1)(106));
F2107: entity F port map(lamdaA => P(2)(107),lamdaB => P(2)(235),lamdaOut => P(1)(107));
F2108: entity F port map(lamdaA => P(2)(108),lamdaB => P(2)(236),lamdaOut => P(1)(108));
F2109: entity F port map(lamdaA => P(2)(109),lamdaB => P(2)(237),lamdaOut => P(1)(109));
F2110: entity F port map(lamdaA => P(2)(110),lamdaB => P(2)(238),lamdaOut => P(1)(110));
F2111: entity F port map(lamdaA => P(2)(111),lamdaB => P(2)(239),lamdaOut => P(1)(111));
F2112: entity F port map(lamdaA => P(2)(112),lamdaB => P(2)(240),lamdaOut => P(1)(112));
F2113: entity F port map(lamdaA => P(2)(113),lamdaB => P(2)(241),lamdaOut => P(1)(113));
F2114: entity F port map(lamdaA => P(2)(114),lamdaB => P(2)(242),lamdaOut => P(1)(114));
F2115: entity F port map(lamdaA => P(2)(115),lamdaB => P(2)(243),lamdaOut => P(1)(115));
F2116: entity F port map(lamdaA => P(2)(116),lamdaB => P(2)(244),lamdaOut => P(1)(116));
F2117: entity F port map(lamdaA => P(2)(117),lamdaB => P(2)(245),lamdaOut => P(1)(117));
F2118: entity F port map(lamdaA => P(2)(118),lamdaB => P(2)(246),lamdaOut => P(1)(118));
F2119: entity F port map(lamdaA => P(2)(119),lamdaB => P(2)(247),lamdaOut => P(1)(119));
F2120: entity F port map(lamdaA => P(2)(120),lamdaB => P(2)(248),lamdaOut => P(1)(120));
F2121: entity F port map(lamdaA => P(2)(121),lamdaB => P(2)(249),lamdaOut => P(1)(121));
F2122: entity F port map(lamdaA => P(2)(122),lamdaB => P(2)(250),lamdaOut => P(1)(122));
F2123: entity F port map(lamdaA => P(2)(123),lamdaB => P(2)(251),lamdaOut => P(1)(123));
F2124: entity F port map(lamdaA => P(2)(124),lamdaB => P(2)(252),lamdaOut => P(1)(124));
F2125: entity F port map(lamdaA => P(2)(125),lamdaB => P(2)(253),lamdaOut => P(1)(125));
F2126: entity F port map(lamdaA => P(2)(126),lamdaB => P(2)(254),lamdaOut => P(1)(126));
F2127: entity F port map(lamdaA => P(2)(127),lamdaB => P(2)(255),lamdaOut => P(1)(127));
G2128: entity G port map(lamdaA => P(2)(0),lamdaB => P(2)(128),s => s(2)(0),lamdaOut => P(1)(128));
G2129: entity G port map(lamdaA => P(2)(1),lamdaB => P(2)(129),s => s(2)(1),lamdaOut => P(1)(129));
G2130: entity G port map(lamdaA => P(2)(2),lamdaB => P(2)(130),s => s(2)(2),lamdaOut => P(1)(130));
G2131: entity G port map(lamdaA => P(2)(3),lamdaB => P(2)(131),s => s(2)(3),lamdaOut => P(1)(131));
G2132: entity G port map(lamdaA => P(2)(4),lamdaB => P(2)(132),s => s(2)(4),lamdaOut => P(1)(132));
G2133: entity G port map(lamdaA => P(2)(5),lamdaB => P(2)(133),s => s(2)(5),lamdaOut => P(1)(133));
G2134: entity G port map(lamdaA => P(2)(6),lamdaB => P(2)(134),s => s(2)(6),lamdaOut => P(1)(134));
G2135: entity G port map(lamdaA => P(2)(7),lamdaB => P(2)(135),s => s(2)(7),lamdaOut => P(1)(135));
G2136: entity G port map(lamdaA => P(2)(8),lamdaB => P(2)(136),s => s(2)(8),lamdaOut => P(1)(136));
G2137: entity G port map(lamdaA => P(2)(9),lamdaB => P(2)(137),s => s(2)(9),lamdaOut => P(1)(137));
G2138: entity G port map(lamdaA => P(2)(10),lamdaB => P(2)(138),s => s(2)(10),lamdaOut => P(1)(138));
G2139: entity G port map(lamdaA => P(2)(11),lamdaB => P(2)(139),s => s(2)(11),lamdaOut => P(1)(139));
G2140: entity G port map(lamdaA => P(2)(12),lamdaB => P(2)(140),s => s(2)(12),lamdaOut => P(1)(140));
G2141: entity G port map(lamdaA => P(2)(13),lamdaB => P(2)(141),s => s(2)(13),lamdaOut => P(1)(141));
G2142: entity G port map(lamdaA => P(2)(14),lamdaB => P(2)(142),s => s(2)(14),lamdaOut => P(1)(142));
G2143: entity G port map(lamdaA => P(2)(15),lamdaB => P(2)(143),s => s(2)(15),lamdaOut => P(1)(143));
G2144: entity G port map(lamdaA => P(2)(16),lamdaB => P(2)(144),s => s(2)(16),lamdaOut => P(1)(144));
G2145: entity G port map(lamdaA => P(2)(17),lamdaB => P(2)(145),s => s(2)(17),lamdaOut => P(1)(145));
G2146: entity G port map(lamdaA => P(2)(18),lamdaB => P(2)(146),s => s(2)(18),lamdaOut => P(1)(146));
G2147: entity G port map(lamdaA => P(2)(19),lamdaB => P(2)(147),s => s(2)(19),lamdaOut => P(1)(147));
G2148: entity G port map(lamdaA => P(2)(20),lamdaB => P(2)(148),s => s(2)(20),lamdaOut => P(1)(148));
G2149: entity G port map(lamdaA => P(2)(21),lamdaB => P(2)(149),s => s(2)(21),lamdaOut => P(1)(149));
G2150: entity G port map(lamdaA => P(2)(22),lamdaB => P(2)(150),s => s(2)(22),lamdaOut => P(1)(150));
G2151: entity G port map(lamdaA => P(2)(23),lamdaB => P(2)(151),s => s(2)(23),lamdaOut => P(1)(151));
G2152: entity G port map(lamdaA => P(2)(24),lamdaB => P(2)(152),s => s(2)(24),lamdaOut => P(1)(152));
G2153: entity G port map(lamdaA => P(2)(25),lamdaB => P(2)(153),s => s(2)(25),lamdaOut => P(1)(153));
G2154: entity G port map(lamdaA => P(2)(26),lamdaB => P(2)(154),s => s(2)(26),lamdaOut => P(1)(154));
G2155: entity G port map(lamdaA => P(2)(27),lamdaB => P(2)(155),s => s(2)(27),lamdaOut => P(1)(155));
G2156: entity G port map(lamdaA => P(2)(28),lamdaB => P(2)(156),s => s(2)(28),lamdaOut => P(1)(156));
G2157: entity G port map(lamdaA => P(2)(29),lamdaB => P(2)(157),s => s(2)(29),lamdaOut => P(1)(157));
G2158: entity G port map(lamdaA => P(2)(30),lamdaB => P(2)(158),s => s(2)(30),lamdaOut => P(1)(158));
G2159: entity G port map(lamdaA => P(2)(31),lamdaB => P(2)(159),s => s(2)(31),lamdaOut => P(1)(159));
G2160: entity G port map(lamdaA => P(2)(32),lamdaB => P(2)(160),s => s(2)(32),lamdaOut => P(1)(160));
G2161: entity G port map(lamdaA => P(2)(33),lamdaB => P(2)(161),s => s(2)(33),lamdaOut => P(1)(161));
G2162: entity G port map(lamdaA => P(2)(34),lamdaB => P(2)(162),s => s(2)(34),lamdaOut => P(1)(162));
G2163: entity G port map(lamdaA => P(2)(35),lamdaB => P(2)(163),s => s(2)(35),lamdaOut => P(1)(163));
G2164: entity G port map(lamdaA => P(2)(36),lamdaB => P(2)(164),s => s(2)(36),lamdaOut => P(1)(164));
G2165: entity G port map(lamdaA => P(2)(37),lamdaB => P(2)(165),s => s(2)(37),lamdaOut => P(1)(165));
G2166: entity G port map(lamdaA => P(2)(38),lamdaB => P(2)(166),s => s(2)(38),lamdaOut => P(1)(166));
G2167: entity G port map(lamdaA => P(2)(39),lamdaB => P(2)(167),s => s(2)(39),lamdaOut => P(1)(167));
G2168: entity G port map(lamdaA => P(2)(40),lamdaB => P(2)(168),s => s(2)(40),lamdaOut => P(1)(168));
G2169: entity G port map(lamdaA => P(2)(41),lamdaB => P(2)(169),s => s(2)(41),lamdaOut => P(1)(169));
G2170: entity G port map(lamdaA => P(2)(42),lamdaB => P(2)(170),s => s(2)(42),lamdaOut => P(1)(170));
G2171: entity G port map(lamdaA => P(2)(43),lamdaB => P(2)(171),s => s(2)(43),lamdaOut => P(1)(171));
G2172: entity G port map(lamdaA => P(2)(44),lamdaB => P(2)(172),s => s(2)(44),lamdaOut => P(1)(172));
G2173: entity G port map(lamdaA => P(2)(45),lamdaB => P(2)(173),s => s(2)(45),lamdaOut => P(1)(173));
G2174: entity G port map(lamdaA => P(2)(46),lamdaB => P(2)(174),s => s(2)(46),lamdaOut => P(1)(174));
G2175: entity G port map(lamdaA => P(2)(47),lamdaB => P(2)(175),s => s(2)(47),lamdaOut => P(1)(175));
G2176: entity G port map(lamdaA => P(2)(48),lamdaB => P(2)(176),s => s(2)(48),lamdaOut => P(1)(176));
G2177: entity G port map(lamdaA => P(2)(49),lamdaB => P(2)(177),s => s(2)(49),lamdaOut => P(1)(177));
G2178: entity G port map(lamdaA => P(2)(50),lamdaB => P(2)(178),s => s(2)(50),lamdaOut => P(1)(178));
G2179: entity G port map(lamdaA => P(2)(51),lamdaB => P(2)(179),s => s(2)(51),lamdaOut => P(1)(179));
G2180: entity G port map(lamdaA => P(2)(52),lamdaB => P(2)(180),s => s(2)(52),lamdaOut => P(1)(180));
G2181: entity G port map(lamdaA => P(2)(53),lamdaB => P(2)(181),s => s(2)(53),lamdaOut => P(1)(181));
G2182: entity G port map(lamdaA => P(2)(54),lamdaB => P(2)(182),s => s(2)(54),lamdaOut => P(1)(182));
G2183: entity G port map(lamdaA => P(2)(55),lamdaB => P(2)(183),s => s(2)(55),lamdaOut => P(1)(183));
G2184: entity G port map(lamdaA => P(2)(56),lamdaB => P(2)(184),s => s(2)(56),lamdaOut => P(1)(184));
G2185: entity G port map(lamdaA => P(2)(57),lamdaB => P(2)(185),s => s(2)(57),lamdaOut => P(1)(185));
G2186: entity G port map(lamdaA => P(2)(58),lamdaB => P(2)(186),s => s(2)(58),lamdaOut => P(1)(186));
G2187: entity G port map(lamdaA => P(2)(59),lamdaB => P(2)(187),s => s(2)(59),lamdaOut => P(1)(187));
G2188: entity G port map(lamdaA => P(2)(60),lamdaB => P(2)(188),s => s(2)(60),lamdaOut => P(1)(188));
G2189: entity G port map(lamdaA => P(2)(61),lamdaB => P(2)(189),s => s(2)(61),lamdaOut => P(1)(189));
G2190: entity G port map(lamdaA => P(2)(62),lamdaB => P(2)(190),s => s(2)(62),lamdaOut => P(1)(190));
G2191: entity G port map(lamdaA => P(2)(63),lamdaB => P(2)(191),s => s(2)(63),lamdaOut => P(1)(191));
G2192: entity G port map(lamdaA => P(2)(64),lamdaB => P(2)(192),s => s(2)(64),lamdaOut => P(1)(192));
G2193: entity G port map(lamdaA => P(2)(65),lamdaB => P(2)(193),s => s(2)(65),lamdaOut => P(1)(193));
G2194: entity G port map(lamdaA => P(2)(66),lamdaB => P(2)(194),s => s(2)(66),lamdaOut => P(1)(194));
G2195: entity G port map(lamdaA => P(2)(67),lamdaB => P(2)(195),s => s(2)(67),lamdaOut => P(1)(195));
G2196: entity G port map(lamdaA => P(2)(68),lamdaB => P(2)(196),s => s(2)(68),lamdaOut => P(1)(196));
G2197: entity G port map(lamdaA => P(2)(69),lamdaB => P(2)(197),s => s(2)(69),lamdaOut => P(1)(197));
G2198: entity G port map(lamdaA => P(2)(70),lamdaB => P(2)(198),s => s(2)(70),lamdaOut => P(1)(198));
G2199: entity G port map(lamdaA => P(2)(71),lamdaB => P(2)(199),s => s(2)(71),lamdaOut => P(1)(199));
G2200: entity G port map(lamdaA => P(2)(72),lamdaB => P(2)(200),s => s(2)(72),lamdaOut => P(1)(200));
G2201: entity G port map(lamdaA => P(2)(73),lamdaB => P(2)(201),s => s(2)(73),lamdaOut => P(1)(201));
G2202: entity G port map(lamdaA => P(2)(74),lamdaB => P(2)(202),s => s(2)(74),lamdaOut => P(1)(202));
G2203: entity G port map(lamdaA => P(2)(75),lamdaB => P(2)(203),s => s(2)(75),lamdaOut => P(1)(203));
G2204: entity G port map(lamdaA => P(2)(76),lamdaB => P(2)(204),s => s(2)(76),lamdaOut => P(1)(204));
G2205: entity G port map(lamdaA => P(2)(77),lamdaB => P(2)(205),s => s(2)(77),lamdaOut => P(1)(205));
G2206: entity G port map(lamdaA => P(2)(78),lamdaB => P(2)(206),s => s(2)(78),lamdaOut => P(1)(206));
G2207: entity G port map(lamdaA => P(2)(79),lamdaB => P(2)(207),s => s(2)(79),lamdaOut => P(1)(207));
G2208: entity G port map(lamdaA => P(2)(80),lamdaB => P(2)(208),s => s(2)(80),lamdaOut => P(1)(208));
G2209: entity G port map(lamdaA => P(2)(81),lamdaB => P(2)(209),s => s(2)(81),lamdaOut => P(1)(209));
G2210: entity G port map(lamdaA => P(2)(82),lamdaB => P(2)(210),s => s(2)(82),lamdaOut => P(1)(210));
G2211: entity G port map(lamdaA => P(2)(83),lamdaB => P(2)(211),s => s(2)(83),lamdaOut => P(1)(211));
G2212: entity G port map(lamdaA => P(2)(84),lamdaB => P(2)(212),s => s(2)(84),lamdaOut => P(1)(212));
G2213: entity G port map(lamdaA => P(2)(85),lamdaB => P(2)(213),s => s(2)(85),lamdaOut => P(1)(213));
G2214: entity G port map(lamdaA => P(2)(86),lamdaB => P(2)(214),s => s(2)(86),lamdaOut => P(1)(214));
G2215: entity G port map(lamdaA => P(2)(87),lamdaB => P(2)(215),s => s(2)(87),lamdaOut => P(1)(215));
G2216: entity G port map(lamdaA => P(2)(88),lamdaB => P(2)(216),s => s(2)(88),lamdaOut => P(1)(216));
G2217: entity G port map(lamdaA => P(2)(89),lamdaB => P(2)(217),s => s(2)(89),lamdaOut => P(1)(217));
G2218: entity G port map(lamdaA => P(2)(90),lamdaB => P(2)(218),s => s(2)(90),lamdaOut => P(1)(218));
G2219: entity G port map(lamdaA => P(2)(91),lamdaB => P(2)(219),s => s(2)(91),lamdaOut => P(1)(219));
G2220: entity G port map(lamdaA => P(2)(92),lamdaB => P(2)(220),s => s(2)(92),lamdaOut => P(1)(220));
G2221: entity G port map(lamdaA => P(2)(93),lamdaB => P(2)(221),s => s(2)(93),lamdaOut => P(1)(221));
G2222: entity G port map(lamdaA => P(2)(94),lamdaB => P(2)(222),s => s(2)(94),lamdaOut => P(1)(222));
G2223: entity G port map(lamdaA => P(2)(95),lamdaB => P(2)(223),s => s(2)(95),lamdaOut => P(1)(223));
G2224: entity G port map(lamdaA => P(2)(96),lamdaB => P(2)(224),s => s(2)(96),lamdaOut => P(1)(224));
G2225: entity G port map(lamdaA => P(2)(97),lamdaB => P(2)(225),s => s(2)(97),lamdaOut => P(1)(225));
G2226: entity G port map(lamdaA => P(2)(98),lamdaB => P(2)(226),s => s(2)(98),lamdaOut => P(1)(226));
G2227: entity G port map(lamdaA => P(2)(99),lamdaB => P(2)(227),s => s(2)(99),lamdaOut => P(1)(227));
G2228: entity G port map(lamdaA => P(2)(100),lamdaB => P(2)(228),s => s(2)(100),lamdaOut => P(1)(228));
G2229: entity G port map(lamdaA => P(2)(101),lamdaB => P(2)(229),s => s(2)(101),lamdaOut => P(1)(229));
G2230: entity G port map(lamdaA => P(2)(102),lamdaB => P(2)(230),s => s(2)(102),lamdaOut => P(1)(230));
G2231: entity G port map(lamdaA => P(2)(103),lamdaB => P(2)(231),s => s(2)(103),lamdaOut => P(1)(231));
G2232: entity G port map(lamdaA => P(2)(104),lamdaB => P(2)(232),s => s(2)(104),lamdaOut => P(1)(232));
G2233: entity G port map(lamdaA => P(2)(105),lamdaB => P(2)(233),s => s(2)(105),lamdaOut => P(1)(233));
G2234: entity G port map(lamdaA => P(2)(106),lamdaB => P(2)(234),s => s(2)(106),lamdaOut => P(1)(234));
G2235: entity G port map(lamdaA => P(2)(107),lamdaB => P(2)(235),s => s(2)(107),lamdaOut => P(1)(235));
G2236: entity G port map(lamdaA => P(2)(108),lamdaB => P(2)(236),s => s(2)(108),lamdaOut => P(1)(236));
G2237: entity G port map(lamdaA => P(2)(109),lamdaB => P(2)(237),s => s(2)(109),lamdaOut => P(1)(237));
G2238: entity G port map(lamdaA => P(2)(110),lamdaB => P(2)(238),s => s(2)(110),lamdaOut => P(1)(238));
G2239: entity G port map(lamdaA => P(2)(111),lamdaB => P(2)(239),s => s(2)(111),lamdaOut => P(1)(239));
G2240: entity G port map(lamdaA => P(2)(112),lamdaB => P(2)(240),s => s(2)(112),lamdaOut => P(1)(240));
G2241: entity G port map(lamdaA => P(2)(113),lamdaB => P(2)(241),s => s(2)(113),lamdaOut => P(1)(241));
G2242: entity G port map(lamdaA => P(2)(114),lamdaB => P(2)(242),s => s(2)(114),lamdaOut => P(1)(242));
G2243: entity G port map(lamdaA => P(2)(115),lamdaB => P(2)(243),s => s(2)(115),lamdaOut => P(1)(243));
G2244: entity G port map(lamdaA => P(2)(116),lamdaB => P(2)(244),s => s(2)(116),lamdaOut => P(1)(244));
G2245: entity G port map(lamdaA => P(2)(117),lamdaB => P(2)(245),s => s(2)(117),lamdaOut => P(1)(245));
G2246: entity G port map(lamdaA => P(2)(118),lamdaB => P(2)(246),s => s(2)(118),lamdaOut => P(1)(246));
G2247: entity G port map(lamdaA => P(2)(119),lamdaB => P(2)(247),s => s(2)(119),lamdaOut => P(1)(247));
G2248: entity G port map(lamdaA => P(2)(120),lamdaB => P(2)(248),s => s(2)(120),lamdaOut => P(1)(248));
G2249: entity G port map(lamdaA => P(2)(121),lamdaB => P(2)(249),s => s(2)(121),lamdaOut => P(1)(249));
G2250: entity G port map(lamdaA => P(2)(122),lamdaB => P(2)(250),s => s(2)(122),lamdaOut => P(1)(250));
G2251: entity G port map(lamdaA => P(2)(123),lamdaB => P(2)(251),s => s(2)(123),lamdaOut => P(1)(251));
G2252: entity G port map(lamdaA => P(2)(124),lamdaB => P(2)(252),s => s(2)(124),lamdaOut => P(1)(252));
G2253: entity G port map(lamdaA => P(2)(125),lamdaB => P(2)(253),s => s(2)(125),lamdaOut => P(1)(253));
G2254: entity G port map(lamdaA => P(2)(126),lamdaB => P(2)(254),s => s(2)(126),lamdaOut => P(1)(254));
G2255: entity G port map(lamdaA => P(2)(127),lamdaB => P(2)(255),s => s(2)(127),lamdaOut => P(1)(255));
F2256: entity F port map(lamdaA => P(2)(256),lamdaB => P(2)(384),lamdaOut => P(1)(256));
F2257: entity F port map(lamdaA => P(2)(257),lamdaB => P(2)(385),lamdaOut => P(1)(257));
F2258: entity F port map(lamdaA => P(2)(258),lamdaB => P(2)(386),lamdaOut => P(1)(258));
F2259: entity F port map(lamdaA => P(2)(259),lamdaB => P(2)(387),lamdaOut => P(1)(259));
F2260: entity F port map(lamdaA => P(2)(260),lamdaB => P(2)(388),lamdaOut => P(1)(260));
F2261: entity F port map(lamdaA => P(2)(261),lamdaB => P(2)(389),lamdaOut => P(1)(261));
F2262: entity F port map(lamdaA => P(2)(262),lamdaB => P(2)(390),lamdaOut => P(1)(262));
F2263: entity F port map(lamdaA => P(2)(263),lamdaB => P(2)(391),lamdaOut => P(1)(263));
F2264: entity F port map(lamdaA => P(2)(264),lamdaB => P(2)(392),lamdaOut => P(1)(264));
F2265: entity F port map(lamdaA => P(2)(265),lamdaB => P(2)(393),lamdaOut => P(1)(265));
F2266: entity F port map(lamdaA => P(2)(266),lamdaB => P(2)(394),lamdaOut => P(1)(266));
F2267: entity F port map(lamdaA => P(2)(267),lamdaB => P(2)(395),lamdaOut => P(1)(267));
F2268: entity F port map(lamdaA => P(2)(268),lamdaB => P(2)(396),lamdaOut => P(1)(268));
F2269: entity F port map(lamdaA => P(2)(269),lamdaB => P(2)(397),lamdaOut => P(1)(269));
F2270: entity F port map(lamdaA => P(2)(270),lamdaB => P(2)(398),lamdaOut => P(1)(270));
F2271: entity F port map(lamdaA => P(2)(271),lamdaB => P(2)(399),lamdaOut => P(1)(271));
F2272: entity F port map(lamdaA => P(2)(272),lamdaB => P(2)(400),lamdaOut => P(1)(272));
F2273: entity F port map(lamdaA => P(2)(273),lamdaB => P(2)(401),lamdaOut => P(1)(273));
F2274: entity F port map(lamdaA => P(2)(274),lamdaB => P(2)(402),lamdaOut => P(1)(274));
F2275: entity F port map(lamdaA => P(2)(275),lamdaB => P(2)(403),lamdaOut => P(1)(275));
F2276: entity F port map(lamdaA => P(2)(276),lamdaB => P(2)(404),lamdaOut => P(1)(276));
F2277: entity F port map(lamdaA => P(2)(277),lamdaB => P(2)(405),lamdaOut => P(1)(277));
F2278: entity F port map(lamdaA => P(2)(278),lamdaB => P(2)(406),lamdaOut => P(1)(278));
F2279: entity F port map(lamdaA => P(2)(279),lamdaB => P(2)(407),lamdaOut => P(1)(279));
F2280: entity F port map(lamdaA => P(2)(280),lamdaB => P(2)(408),lamdaOut => P(1)(280));
F2281: entity F port map(lamdaA => P(2)(281),lamdaB => P(2)(409),lamdaOut => P(1)(281));
F2282: entity F port map(lamdaA => P(2)(282),lamdaB => P(2)(410),lamdaOut => P(1)(282));
F2283: entity F port map(lamdaA => P(2)(283),lamdaB => P(2)(411),lamdaOut => P(1)(283));
F2284: entity F port map(lamdaA => P(2)(284),lamdaB => P(2)(412),lamdaOut => P(1)(284));
F2285: entity F port map(lamdaA => P(2)(285),lamdaB => P(2)(413),lamdaOut => P(1)(285));
F2286: entity F port map(lamdaA => P(2)(286),lamdaB => P(2)(414),lamdaOut => P(1)(286));
F2287: entity F port map(lamdaA => P(2)(287),lamdaB => P(2)(415),lamdaOut => P(1)(287));
F2288: entity F port map(lamdaA => P(2)(288),lamdaB => P(2)(416),lamdaOut => P(1)(288));
F2289: entity F port map(lamdaA => P(2)(289),lamdaB => P(2)(417),lamdaOut => P(1)(289));
F2290: entity F port map(lamdaA => P(2)(290),lamdaB => P(2)(418),lamdaOut => P(1)(290));
F2291: entity F port map(lamdaA => P(2)(291),lamdaB => P(2)(419),lamdaOut => P(1)(291));
F2292: entity F port map(lamdaA => P(2)(292),lamdaB => P(2)(420),lamdaOut => P(1)(292));
F2293: entity F port map(lamdaA => P(2)(293),lamdaB => P(2)(421),lamdaOut => P(1)(293));
F2294: entity F port map(lamdaA => P(2)(294),lamdaB => P(2)(422),lamdaOut => P(1)(294));
F2295: entity F port map(lamdaA => P(2)(295),lamdaB => P(2)(423),lamdaOut => P(1)(295));
F2296: entity F port map(lamdaA => P(2)(296),lamdaB => P(2)(424),lamdaOut => P(1)(296));
F2297: entity F port map(lamdaA => P(2)(297),lamdaB => P(2)(425),lamdaOut => P(1)(297));
F2298: entity F port map(lamdaA => P(2)(298),lamdaB => P(2)(426),lamdaOut => P(1)(298));
F2299: entity F port map(lamdaA => P(2)(299),lamdaB => P(2)(427),lamdaOut => P(1)(299));
F2300: entity F port map(lamdaA => P(2)(300),lamdaB => P(2)(428),lamdaOut => P(1)(300));
F2301: entity F port map(lamdaA => P(2)(301),lamdaB => P(2)(429),lamdaOut => P(1)(301));
F2302: entity F port map(lamdaA => P(2)(302),lamdaB => P(2)(430),lamdaOut => P(1)(302));
F2303: entity F port map(lamdaA => P(2)(303),lamdaB => P(2)(431),lamdaOut => P(1)(303));
F2304: entity F port map(lamdaA => P(2)(304),lamdaB => P(2)(432),lamdaOut => P(1)(304));
F2305: entity F port map(lamdaA => P(2)(305),lamdaB => P(2)(433),lamdaOut => P(1)(305));
F2306: entity F port map(lamdaA => P(2)(306),lamdaB => P(2)(434),lamdaOut => P(1)(306));
F2307: entity F port map(lamdaA => P(2)(307),lamdaB => P(2)(435),lamdaOut => P(1)(307));
F2308: entity F port map(lamdaA => P(2)(308),lamdaB => P(2)(436),lamdaOut => P(1)(308));
F2309: entity F port map(lamdaA => P(2)(309),lamdaB => P(2)(437),lamdaOut => P(1)(309));
F2310: entity F port map(lamdaA => P(2)(310),lamdaB => P(2)(438),lamdaOut => P(1)(310));
F2311: entity F port map(lamdaA => P(2)(311),lamdaB => P(2)(439),lamdaOut => P(1)(311));
F2312: entity F port map(lamdaA => P(2)(312),lamdaB => P(2)(440),lamdaOut => P(1)(312));
F2313: entity F port map(lamdaA => P(2)(313),lamdaB => P(2)(441),lamdaOut => P(1)(313));
F2314: entity F port map(lamdaA => P(2)(314),lamdaB => P(2)(442),lamdaOut => P(1)(314));
F2315: entity F port map(lamdaA => P(2)(315),lamdaB => P(2)(443),lamdaOut => P(1)(315));
F2316: entity F port map(lamdaA => P(2)(316),lamdaB => P(2)(444),lamdaOut => P(1)(316));
F2317: entity F port map(lamdaA => P(2)(317),lamdaB => P(2)(445),lamdaOut => P(1)(317));
F2318: entity F port map(lamdaA => P(2)(318),lamdaB => P(2)(446),lamdaOut => P(1)(318));
F2319: entity F port map(lamdaA => P(2)(319),lamdaB => P(2)(447),lamdaOut => P(1)(319));
F2320: entity F port map(lamdaA => P(2)(320),lamdaB => P(2)(448),lamdaOut => P(1)(320));
F2321: entity F port map(lamdaA => P(2)(321),lamdaB => P(2)(449),lamdaOut => P(1)(321));
F2322: entity F port map(lamdaA => P(2)(322),lamdaB => P(2)(450),lamdaOut => P(1)(322));
F2323: entity F port map(lamdaA => P(2)(323),lamdaB => P(2)(451),lamdaOut => P(1)(323));
F2324: entity F port map(lamdaA => P(2)(324),lamdaB => P(2)(452),lamdaOut => P(1)(324));
F2325: entity F port map(lamdaA => P(2)(325),lamdaB => P(2)(453),lamdaOut => P(1)(325));
F2326: entity F port map(lamdaA => P(2)(326),lamdaB => P(2)(454),lamdaOut => P(1)(326));
F2327: entity F port map(lamdaA => P(2)(327),lamdaB => P(2)(455),lamdaOut => P(1)(327));
F2328: entity F port map(lamdaA => P(2)(328),lamdaB => P(2)(456),lamdaOut => P(1)(328));
F2329: entity F port map(lamdaA => P(2)(329),lamdaB => P(2)(457),lamdaOut => P(1)(329));
F2330: entity F port map(lamdaA => P(2)(330),lamdaB => P(2)(458),lamdaOut => P(1)(330));
F2331: entity F port map(lamdaA => P(2)(331),lamdaB => P(2)(459),lamdaOut => P(1)(331));
F2332: entity F port map(lamdaA => P(2)(332),lamdaB => P(2)(460),lamdaOut => P(1)(332));
F2333: entity F port map(lamdaA => P(2)(333),lamdaB => P(2)(461),lamdaOut => P(1)(333));
F2334: entity F port map(lamdaA => P(2)(334),lamdaB => P(2)(462),lamdaOut => P(1)(334));
F2335: entity F port map(lamdaA => P(2)(335),lamdaB => P(2)(463),lamdaOut => P(1)(335));
F2336: entity F port map(lamdaA => P(2)(336),lamdaB => P(2)(464),lamdaOut => P(1)(336));
F2337: entity F port map(lamdaA => P(2)(337),lamdaB => P(2)(465),lamdaOut => P(1)(337));
F2338: entity F port map(lamdaA => P(2)(338),lamdaB => P(2)(466),lamdaOut => P(1)(338));
F2339: entity F port map(lamdaA => P(2)(339),lamdaB => P(2)(467),lamdaOut => P(1)(339));
F2340: entity F port map(lamdaA => P(2)(340),lamdaB => P(2)(468),lamdaOut => P(1)(340));
F2341: entity F port map(lamdaA => P(2)(341),lamdaB => P(2)(469),lamdaOut => P(1)(341));
F2342: entity F port map(lamdaA => P(2)(342),lamdaB => P(2)(470),lamdaOut => P(1)(342));
F2343: entity F port map(lamdaA => P(2)(343),lamdaB => P(2)(471),lamdaOut => P(1)(343));
F2344: entity F port map(lamdaA => P(2)(344),lamdaB => P(2)(472),lamdaOut => P(1)(344));
F2345: entity F port map(lamdaA => P(2)(345),lamdaB => P(2)(473),lamdaOut => P(1)(345));
F2346: entity F port map(lamdaA => P(2)(346),lamdaB => P(2)(474),lamdaOut => P(1)(346));
F2347: entity F port map(lamdaA => P(2)(347),lamdaB => P(2)(475),lamdaOut => P(1)(347));
F2348: entity F port map(lamdaA => P(2)(348),lamdaB => P(2)(476),lamdaOut => P(1)(348));
F2349: entity F port map(lamdaA => P(2)(349),lamdaB => P(2)(477),lamdaOut => P(1)(349));
F2350: entity F port map(lamdaA => P(2)(350),lamdaB => P(2)(478),lamdaOut => P(1)(350));
F2351: entity F port map(lamdaA => P(2)(351),lamdaB => P(2)(479),lamdaOut => P(1)(351));
F2352: entity F port map(lamdaA => P(2)(352),lamdaB => P(2)(480),lamdaOut => P(1)(352));
F2353: entity F port map(lamdaA => P(2)(353),lamdaB => P(2)(481),lamdaOut => P(1)(353));
F2354: entity F port map(lamdaA => P(2)(354),lamdaB => P(2)(482),lamdaOut => P(1)(354));
F2355: entity F port map(lamdaA => P(2)(355),lamdaB => P(2)(483),lamdaOut => P(1)(355));
F2356: entity F port map(lamdaA => P(2)(356),lamdaB => P(2)(484),lamdaOut => P(1)(356));
F2357: entity F port map(lamdaA => P(2)(357),lamdaB => P(2)(485),lamdaOut => P(1)(357));
F2358: entity F port map(lamdaA => P(2)(358),lamdaB => P(2)(486),lamdaOut => P(1)(358));
F2359: entity F port map(lamdaA => P(2)(359),lamdaB => P(2)(487),lamdaOut => P(1)(359));
F2360: entity F port map(lamdaA => P(2)(360),lamdaB => P(2)(488),lamdaOut => P(1)(360));
F2361: entity F port map(lamdaA => P(2)(361),lamdaB => P(2)(489),lamdaOut => P(1)(361));
F2362: entity F port map(lamdaA => P(2)(362),lamdaB => P(2)(490),lamdaOut => P(1)(362));
F2363: entity F port map(lamdaA => P(2)(363),lamdaB => P(2)(491),lamdaOut => P(1)(363));
F2364: entity F port map(lamdaA => P(2)(364),lamdaB => P(2)(492),lamdaOut => P(1)(364));
F2365: entity F port map(lamdaA => P(2)(365),lamdaB => P(2)(493),lamdaOut => P(1)(365));
F2366: entity F port map(lamdaA => P(2)(366),lamdaB => P(2)(494),lamdaOut => P(1)(366));
F2367: entity F port map(lamdaA => P(2)(367),lamdaB => P(2)(495),lamdaOut => P(1)(367));
F2368: entity F port map(lamdaA => P(2)(368),lamdaB => P(2)(496),lamdaOut => P(1)(368));
F2369: entity F port map(lamdaA => P(2)(369),lamdaB => P(2)(497),lamdaOut => P(1)(369));
F2370: entity F port map(lamdaA => P(2)(370),lamdaB => P(2)(498),lamdaOut => P(1)(370));
F2371: entity F port map(lamdaA => P(2)(371),lamdaB => P(2)(499),lamdaOut => P(1)(371));
F2372: entity F port map(lamdaA => P(2)(372),lamdaB => P(2)(500),lamdaOut => P(1)(372));
F2373: entity F port map(lamdaA => P(2)(373),lamdaB => P(2)(501),lamdaOut => P(1)(373));
F2374: entity F port map(lamdaA => P(2)(374),lamdaB => P(2)(502),lamdaOut => P(1)(374));
F2375: entity F port map(lamdaA => P(2)(375),lamdaB => P(2)(503),lamdaOut => P(1)(375));
F2376: entity F port map(lamdaA => P(2)(376),lamdaB => P(2)(504),lamdaOut => P(1)(376));
F2377: entity F port map(lamdaA => P(2)(377),lamdaB => P(2)(505),lamdaOut => P(1)(377));
F2378: entity F port map(lamdaA => P(2)(378),lamdaB => P(2)(506),lamdaOut => P(1)(378));
F2379: entity F port map(lamdaA => P(2)(379),lamdaB => P(2)(507),lamdaOut => P(1)(379));
F2380: entity F port map(lamdaA => P(2)(380),lamdaB => P(2)(508),lamdaOut => P(1)(380));
F2381: entity F port map(lamdaA => P(2)(381),lamdaB => P(2)(509),lamdaOut => P(1)(381));
F2382: entity F port map(lamdaA => P(2)(382),lamdaB => P(2)(510),lamdaOut => P(1)(382));
F2383: entity F port map(lamdaA => P(2)(383),lamdaB => P(2)(511),lamdaOut => P(1)(383));
G2384: entity G port map(lamdaA => P(2)(256),lamdaB => P(2)(384),s => s(2)(128),lamdaOut => P(1)(384));
G2385: entity G port map(lamdaA => P(2)(257),lamdaB => P(2)(385),s => s(2)(129),lamdaOut => P(1)(385));
G2386: entity G port map(lamdaA => P(2)(258),lamdaB => P(2)(386),s => s(2)(130),lamdaOut => P(1)(386));
G2387: entity G port map(lamdaA => P(2)(259),lamdaB => P(2)(387),s => s(2)(131),lamdaOut => P(1)(387));
G2388: entity G port map(lamdaA => P(2)(260),lamdaB => P(2)(388),s => s(2)(132),lamdaOut => P(1)(388));
G2389: entity G port map(lamdaA => P(2)(261),lamdaB => P(2)(389),s => s(2)(133),lamdaOut => P(1)(389));
G2390: entity G port map(lamdaA => P(2)(262),lamdaB => P(2)(390),s => s(2)(134),lamdaOut => P(1)(390));
G2391: entity G port map(lamdaA => P(2)(263),lamdaB => P(2)(391),s => s(2)(135),lamdaOut => P(1)(391));
G2392: entity G port map(lamdaA => P(2)(264),lamdaB => P(2)(392),s => s(2)(136),lamdaOut => P(1)(392));
G2393: entity G port map(lamdaA => P(2)(265),lamdaB => P(2)(393),s => s(2)(137),lamdaOut => P(1)(393));
G2394: entity G port map(lamdaA => P(2)(266),lamdaB => P(2)(394),s => s(2)(138),lamdaOut => P(1)(394));
G2395: entity G port map(lamdaA => P(2)(267),lamdaB => P(2)(395),s => s(2)(139),lamdaOut => P(1)(395));
G2396: entity G port map(lamdaA => P(2)(268),lamdaB => P(2)(396),s => s(2)(140),lamdaOut => P(1)(396));
G2397: entity G port map(lamdaA => P(2)(269),lamdaB => P(2)(397),s => s(2)(141),lamdaOut => P(1)(397));
G2398: entity G port map(lamdaA => P(2)(270),lamdaB => P(2)(398),s => s(2)(142),lamdaOut => P(1)(398));
G2399: entity G port map(lamdaA => P(2)(271),lamdaB => P(2)(399),s => s(2)(143),lamdaOut => P(1)(399));
G2400: entity G port map(lamdaA => P(2)(272),lamdaB => P(2)(400),s => s(2)(144),lamdaOut => P(1)(400));
G2401: entity G port map(lamdaA => P(2)(273),lamdaB => P(2)(401),s => s(2)(145),lamdaOut => P(1)(401));
G2402: entity G port map(lamdaA => P(2)(274),lamdaB => P(2)(402),s => s(2)(146),lamdaOut => P(1)(402));
G2403: entity G port map(lamdaA => P(2)(275),lamdaB => P(2)(403),s => s(2)(147),lamdaOut => P(1)(403));
G2404: entity G port map(lamdaA => P(2)(276),lamdaB => P(2)(404),s => s(2)(148),lamdaOut => P(1)(404));
G2405: entity G port map(lamdaA => P(2)(277),lamdaB => P(2)(405),s => s(2)(149),lamdaOut => P(1)(405));
G2406: entity G port map(lamdaA => P(2)(278),lamdaB => P(2)(406),s => s(2)(150),lamdaOut => P(1)(406));
G2407: entity G port map(lamdaA => P(2)(279),lamdaB => P(2)(407),s => s(2)(151),lamdaOut => P(1)(407));
G2408: entity G port map(lamdaA => P(2)(280),lamdaB => P(2)(408),s => s(2)(152),lamdaOut => P(1)(408));
G2409: entity G port map(lamdaA => P(2)(281),lamdaB => P(2)(409),s => s(2)(153),lamdaOut => P(1)(409));
G2410: entity G port map(lamdaA => P(2)(282),lamdaB => P(2)(410),s => s(2)(154),lamdaOut => P(1)(410));
G2411: entity G port map(lamdaA => P(2)(283),lamdaB => P(2)(411),s => s(2)(155),lamdaOut => P(1)(411));
G2412: entity G port map(lamdaA => P(2)(284),lamdaB => P(2)(412),s => s(2)(156),lamdaOut => P(1)(412));
G2413: entity G port map(lamdaA => P(2)(285),lamdaB => P(2)(413),s => s(2)(157),lamdaOut => P(1)(413));
G2414: entity G port map(lamdaA => P(2)(286),lamdaB => P(2)(414),s => s(2)(158),lamdaOut => P(1)(414));
G2415: entity G port map(lamdaA => P(2)(287),lamdaB => P(2)(415),s => s(2)(159),lamdaOut => P(1)(415));
G2416: entity G port map(lamdaA => P(2)(288),lamdaB => P(2)(416),s => s(2)(160),lamdaOut => P(1)(416));
G2417: entity G port map(lamdaA => P(2)(289),lamdaB => P(2)(417),s => s(2)(161),lamdaOut => P(1)(417));
G2418: entity G port map(lamdaA => P(2)(290),lamdaB => P(2)(418),s => s(2)(162),lamdaOut => P(1)(418));
G2419: entity G port map(lamdaA => P(2)(291),lamdaB => P(2)(419),s => s(2)(163),lamdaOut => P(1)(419));
G2420: entity G port map(lamdaA => P(2)(292),lamdaB => P(2)(420),s => s(2)(164),lamdaOut => P(1)(420));
G2421: entity G port map(lamdaA => P(2)(293),lamdaB => P(2)(421),s => s(2)(165),lamdaOut => P(1)(421));
G2422: entity G port map(lamdaA => P(2)(294),lamdaB => P(2)(422),s => s(2)(166),lamdaOut => P(1)(422));
G2423: entity G port map(lamdaA => P(2)(295),lamdaB => P(2)(423),s => s(2)(167),lamdaOut => P(1)(423));
G2424: entity G port map(lamdaA => P(2)(296),lamdaB => P(2)(424),s => s(2)(168),lamdaOut => P(1)(424));
G2425: entity G port map(lamdaA => P(2)(297),lamdaB => P(2)(425),s => s(2)(169),lamdaOut => P(1)(425));
G2426: entity G port map(lamdaA => P(2)(298),lamdaB => P(2)(426),s => s(2)(170),lamdaOut => P(1)(426));
G2427: entity G port map(lamdaA => P(2)(299),lamdaB => P(2)(427),s => s(2)(171),lamdaOut => P(1)(427));
G2428: entity G port map(lamdaA => P(2)(300),lamdaB => P(2)(428),s => s(2)(172),lamdaOut => P(1)(428));
G2429: entity G port map(lamdaA => P(2)(301),lamdaB => P(2)(429),s => s(2)(173),lamdaOut => P(1)(429));
G2430: entity G port map(lamdaA => P(2)(302),lamdaB => P(2)(430),s => s(2)(174),lamdaOut => P(1)(430));
G2431: entity G port map(lamdaA => P(2)(303),lamdaB => P(2)(431),s => s(2)(175),lamdaOut => P(1)(431));
G2432: entity G port map(lamdaA => P(2)(304),lamdaB => P(2)(432),s => s(2)(176),lamdaOut => P(1)(432));
G2433: entity G port map(lamdaA => P(2)(305),lamdaB => P(2)(433),s => s(2)(177),lamdaOut => P(1)(433));
G2434: entity G port map(lamdaA => P(2)(306),lamdaB => P(2)(434),s => s(2)(178),lamdaOut => P(1)(434));
G2435: entity G port map(lamdaA => P(2)(307),lamdaB => P(2)(435),s => s(2)(179),lamdaOut => P(1)(435));
G2436: entity G port map(lamdaA => P(2)(308),lamdaB => P(2)(436),s => s(2)(180),lamdaOut => P(1)(436));
G2437: entity G port map(lamdaA => P(2)(309),lamdaB => P(2)(437),s => s(2)(181),lamdaOut => P(1)(437));
G2438: entity G port map(lamdaA => P(2)(310),lamdaB => P(2)(438),s => s(2)(182),lamdaOut => P(1)(438));
G2439: entity G port map(lamdaA => P(2)(311),lamdaB => P(2)(439),s => s(2)(183),lamdaOut => P(1)(439));
G2440: entity G port map(lamdaA => P(2)(312),lamdaB => P(2)(440),s => s(2)(184),lamdaOut => P(1)(440));
G2441: entity G port map(lamdaA => P(2)(313),lamdaB => P(2)(441),s => s(2)(185),lamdaOut => P(1)(441));
G2442: entity G port map(lamdaA => P(2)(314),lamdaB => P(2)(442),s => s(2)(186),lamdaOut => P(1)(442));
G2443: entity G port map(lamdaA => P(2)(315),lamdaB => P(2)(443),s => s(2)(187),lamdaOut => P(1)(443));
G2444: entity G port map(lamdaA => P(2)(316),lamdaB => P(2)(444),s => s(2)(188),lamdaOut => P(1)(444));
G2445: entity G port map(lamdaA => P(2)(317),lamdaB => P(2)(445),s => s(2)(189),lamdaOut => P(1)(445));
G2446: entity G port map(lamdaA => P(2)(318),lamdaB => P(2)(446),s => s(2)(190),lamdaOut => P(1)(446));
G2447: entity G port map(lamdaA => P(2)(319),lamdaB => P(2)(447),s => s(2)(191),lamdaOut => P(1)(447));
G2448: entity G port map(lamdaA => P(2)(320),lamdaB => P(2)(448),s => s(2)(192),lamdaOut => P(1)(448));
G2449: entity G port map(lamdaA => P(2)(321),lamdaB => P(2)(449),s => s(2)(193),lamdaOut => P(1)(449));
G2450: entity G port map(lamdaA => P(2)(322),lamdaB => P(2)(450),s => s(2)(194),lamdaOut => P(1)(450));
G2451: entity G port map(lamdaA => P(2)(323),lamdaB => P(2)(451),s => s(2)(195),lamdaOut => P(1)(451));
G2452: entity G port map(lamdaA => P(2)(324),lamdaB => P(2)(452),s => s(2)(196),lamdaOut => P(1)(452));
G2453: entity G port map(lamdaA => P(2)(325),lamdaB => P(2)(453),s => s(2)(197),lamdaOut => P(1)(453));
G2454: entity G port map(lamdaA => P(2)(326),lamdaB => P(2)(454),s => s(2)(198),lamdaOut => P(1)(454));
G2455: entity G port map(lamdaA => P(2)(327),lamdaB => P(2)(455),s => s(2)(199),lamdaOut => P(1)(455));
G2456: entity G port map(lamdaA => P(2)(328),lamdaB => P(2)(456),s => s(2)(200),lamdaOut => P(1)(456));
G2457: entity G port map(lamdaA => P(2)(329),lamdaB => P(2)(457),s => s(2)(201),lamdaOut => P(1)(457));
G2458: entity G port map(lamdaA => P(2)(330),lamdaB => P(2)(458),s => s(2)(202),lamdaOut => P(1)(458));
G2459: entity G port map(lamdaA => P(2)(331),lamdaB => P(2)(459),s => s(2)(203),lamdaOut => P(1)(459));
G2460: entity G port map(lamdaA => P(2)(332),lamdaB => P(2)(460),s => s(2)(204),lamdaOut => P(1)(460));
G2461: entity G port map(lamdaA => P(2)(333),lamdaB => P(2)(461),s => s(2)(205),lamdaOut => P(1)(461));
G2462: entity G port map(lamdaA => P(2)(334),lamdaB => P(2)(462),s => s(2)(206),lamdaOut => P(1)(462));
G2463: entity G port map(lamdaA => P(2)(335),lamdaB => P(2)(463),s => s(2)(207),lamdaOut => P(1)(463));
G2464: entity G port map(lamdaA => P(2)(336),lamdaB => P(2)(464),s => s(2)(208),lamdaOut => P(1)(464));
G2465: entity G port map(lamdaA => P(2)(337),lamdaB => P(2)(465),s => s(2)(209),lamdaOut => P(1)(465));
G2466: entity G port map(lamdaA => P(2)(338),lamdaB => P(2)(466),s => s(2)(210),lamdaOut => P(1)(466));
G2467: entity G port map(lamdaA => P(2)(339),lamdaB => P(2)(467),s => s(2)(211),lamdaOut => P(1)(467));
G2468: entity G port map(lamdaA => P(2)(340),lamdaB => P(2)(468),s => s(2)(212),lamdaOut => P(1)(468));
G2469: entity G port map(lamdaA => P(2)(341),lamdaB => P(2)(469),s => s(2)(213),lamdaOut => P(1)(469));
G2470: entity G port map(lamdaA => P(2)(342),lamdaB => P(2)(470),s => s(2)(214),lamdaOut => P(1)(470));
G2471: entity G port map(lamdaA => P(2)(343),lamdaB => P(2)(471),s => s(2)(215),lamdaOut => P(1)(471));
G2472: entity G port map(lamdaA => P(2)(344),lamdaB => P(2)(472),s => s(2)(216),lamdaOut => P(1)(472));
G2473: entity G port map(lamdaA => P(2)(345),lamdaB => P(2)(473),s => s(2)(217),lamdaOut => P(1)(473));
G2474: entity G port map(lamdaA => P(2)(346),lamdaB => P(2)(474),s => s(2)(218),lamdaOut => P(1)(474));
G2475: entity G port map(lamdaA => P(2)(347),lamdaB => P(2)(475),s => s(2)(219),lamdaOut => P(1)(475));
G2476: entity G port map(lamdaA => P(2)(348),lamdaB => P(2)(476),s => s(2)(220),lamdaOut => P(1)(476));
G2477: entity G port map(lamdaA => P(2)(349),lamdaB => P(2)(477),s => s(2)(221),lamdaOut => P(1)(477));
G2478: entity G port map(lamdaA => P(2)(350),lamdaB => P(2)(478),s => s(2)(222),lamdaOut => P(1)(478));
G2479: entity G port map(lamdaA => P(2)(351),lamdaB => P(2)(479),s => s(2)(223),lamdaOut => P(1)(479));
G2480: entity G port map(lamdaA => P(2)(352),lamdaB => P(2)(480),s => s(2)(224),lamdaOut => P(1)(480));
G2481: entity G port map(lamdaA => P(2)(353),lamdaB => P(2)(481),s => s(2)(225),lamdaOut => P(1)(481));
G2482: entity G port map(lamdaA => P(2)(354),lamdaB => P(2)(482),s => s(2)(226),lamdaOut => P(1)(482));
G2483: entity G port map(lamdaA => P(2)(355),lamdaB => P(2)(483),s => s(2)(227),lamdaOut => P(1)(483));
G2484: entity G port map(lamdaA => P(2)(356),lamdaB => P(2)(484),s => s(2)(228),lamdaOut => P(1)(484));
G2485: entity G port map(lamdaA => P(2)(357),lamdaB => P(2)(485),s => s(2)(229),lamdaOut => P(1)(485));
G2486: entity G port map(lamdaA => P(2)(358),lamdaB => P(2)(486),s => s(2)(230),lamdaOut => P(1)(486));
G2487: entity G port map(lamdaA => P(2)(359),lamdaB => P(2)(487),s => s(2)(231),lamdaOut => P(1)(487));
G2488: entity G port map(lamdaA => P(2)(360),lamdaB => P(2)(488),s => s(2)(232),lamdaOut => P(1)(488));
G2489: entity G port map(lamdaA => P(2)(361),lamdaB => P(2)(489),s => s(2)(233),lamdaOut => P(1)(489));
G2490: entity G port map(lamdaA => P(2)(362),lamdaB => P(2)(490),s => s(2)(234),lamdaOut => P(1)(490));
G2491: entity G port map(lamdaA => P(2)(363),lamdaB => P(2)(491),s => s(2)(235),lamdaOut => P(1)(491));
G2492: entity G port map(lamdaA => P(2)(364),lamdaB => P(2)(492),s => s(2)(236),lamdaOut => P(1)(492));
G2493: entity G port map(lamdaA => P(2)(365),lamdaB => P(2)(493),s => s(2)(237),lamdaOut => P(1)(493));
G2494: entity G port map(lamdaA => P(2)(366),lamdaB => P(2)(494),s => s(2)(238),lamdaOut => P(1)(494));
G2495: entity G port map(lamdaA => P(2)(367),lamdaB => P(2)(495),s => s(2)(239),lamdaOut => P(1)(495));
G2496: entity G port map(lamdaA => P(2)(368),lamdaB => P(2)(496),s => s(2)(240),lamdaOut => P(1)(496));
G2497: entity G port map(lamdaA => P(2)(369),lamdaB => P(2)(497),s => s(2)(241),lamdaOut => P(1)(497));
G2498: entity G port map(lamdaA => P(2)(370),lamdaB => P(2)(498),s => s(2)(242),lamdaOut => P(1)(498));
G2499: entity G port map(lamdaA => P(2)(371),lamdaB => P(2)(499),s => s(2)(243),lamdaOut => P(1)(499));
G2500: entity G port map(lamdaA => P(2)(372),lamdaB => P(2)(500),s => s(2)(244),lamdaOut => P(1)(500));
G2501: entity G port map(lamdaA => P(2)(373),lamdaB => P(2)(501),s => s(2)(245),lamdaOut => P(1)(501));
G2502: entity G port map(lamdaA => P(2)(374),lamdaB => P(2)(502),s => s(2)(246),lamdaOut => P(1)(502));
G2503: entity G port map(lamdaA => P(2)(375),lamdaB => P(2)(503),s => s(2)(247),lamdaOut => P(1)(503));
G2504: entity G port map(lamdaA => P(2)(376),lamdaB => P(2)(504),s => s(2)(248),lamdaOut => P(1)(504));
G2505: entity G port map(lamdaA => P(2)(377),lamdaB => P(2)(505),s => s(2)(249),lamdaOut => P(1)(505));
G2506: entity G port map(lamdaA => P(2)(378),lamdaB => P(2)(506),s => s(2)(250),lamdaOut => P(1)(506));
G2507: entity G port map(lamdaA => P(2)(379),lamdaB => P(2)(507),s => s(2)(251),lamdaOut => P(1)(507));
G2508: entity G port map(lamdaA => P(2)(380),lamdaB => P(2)(508),s => s(2)(252),lamdaOut => P(1)(508));
G2509: entity G port map(lamdaA => P(2)(381),lamdaB => P(2)(509),s => s(2)(253),lamdaOut => P(1)(509));
G2510: entity G port map(lamdaA => P(2)(382),lamdaB => P(2)(510),s => s(2)(254),lamdaOut => P(1)(510));
G2511: entity G port map(lamdaA => P(2)(383),lamdaB => P(2)(511),s => s(2)(255),lamdaOut => P(1)(511));
-- STAGE 1
F10: entity F port map(lamdaA => P(1)(0),lamdaB => P(1)(256),lamdaOut => P(0)(0));
F11: entity F port map(lamdaA => P(1)(1),lamdaB => P(1)(257),lamdaOut => P(0)(1));
F12: entity F port map(lamdaA => P(1)(2),lamdaB => P(1)(258),lamdaOut => P(0)(2));
F13: entity F port map(lamdaA => P(1)(3),lamdaB => P(1)(259),lamdaOut => P(0)(3));
F14: entity F port map(lamdaA => P(1)(4),lamdaB => P(1)(260),lamdaOut => P(0)(4));
F15: entity F port map(lamdaA => P(1)(5),lamdaB => P(1)(261),lamdaOut => P(0)(5));
F16: entity F port map(lamdaA => P(1)(6),lamdaB => P(1)(262),lamdaOut => P(0)(6));
F17: entity F port map(lamdaA => P(1)(7),lamdaB => P(1)(263),lamdaOut => P(0)(7));
F18: entity F port map(lamdaA => P(1)(8),lamdaB => P(1)(264),lamdaOut => P(0)(8));
F19: entity F port map(lamdaA => P(1)(9),lamdaB => P(1)(265),lamdaOut => P(0)(9));
F110: entity F port map(lamdaA => P(1)(10),lamdaB => P(1)(266),lamdaOut => P(0)(10));
F111: entity F port map(lamdaA => P(1)(11),lamdaB => P(1)(267),lamdaOut => P(0)(11));
F112: entity F port map(lamdaA => P(1)(12),lamdaB => P(1)(268),lamdaOut => P(0)(12));
F113: entity F port map(lamdaA => P(1)(13),lamdaB => P(1)(269),lamdaOut => P(0)(13));
F114: entity F port map(lamdaA => P(1)(14),lamdaB => P(1)(270),lamdaOut => P(0)(14));
F115: entity F port map(lamdaA => P(1)(15),lamdaB => P(1)(271),lamdaOut => P(0)(15));
F116: entity F port map(lamdaA => P(1)(16),lamdaB => P(1)(272),lamdaOut => P(0)(16));
F117: entity F port map(lamdaA => P(1)(17),lamdaB => P(1)(273),lamdaOut => P(0)(17));
F118: entity F port map(lamdaA => P(1)(18),lamdaB => P(1)(274),lamdaOut => P(0)(18));
F119: entity F port map(lamdaA => P(1)(19),lamdaB => P(1)(275),lamdaOut => P(0)(19));
F120: entity F port map(lamdaA => P(1)(20),lamdaB => P(1)(276),lamdaOut => P(0)(20));
F121: entity F port map(lamdaA => P(1)(21),lamdaB => P(1)(277),lamdaOut => P(0)(21));
F122: entity F port map(lamdaA => P(1)(22),lamdaB => P(1)(278),lamdaOut => P(0)(22));
F123: entity F port map(lamdaA => P(1)(23),lamdaB => P(1)(279),lamdaOut => P(0)(23));
F124: entity F port map(lamdaA => P(1)(24),lamdaB => P(1)(280),lamdaOut => P(0)(24));
F125: entity F port map(lamdaA => P(1)(25),lamdaB => P(1)(281),lamdaOut => P(0)(25));
F126: entity F port map(lamdaA => P(1)(26),lamdaB => P(1)(282),lamdaOut => P(0)(26));
F127: entity F port map(lamdaA => P(1)(27),lamdaB => P(1)(283),lamdaOut => P(0)(27));
F128: entity F port map(lamdaA => P(1)(28),lamdaB => P(1)(284),lamdaOut => P(0)(28));
F129: entity F port map(lamdaA => P(1)(29),lamdaB => P(1)(285),lamdaOut => P(0)(29));
F130: entity F port map(lamdaA => P(1)(30),lamdaB => P(1)(286),lamdaOut => P(0)(30));
F131: entity F port map(lamdaA => P(1)(31),lamdaB => P(1)(287),lamdaOut => P(0)(31));
F132: entity F port map(lamdaA => P(1)(32),lamdaB => P(1)(288),lamdaOut => P(0)(32));
F133: entity F port map(lamdaA => P(1)(33),lamdaB => P(1)(289),lamdaOut => P(0)(33));
F134: entity F port map(lamdaA => P(1)(34),lamdaB => P(1)(290),lamdaOut => P(0)(34));
F135: entity F port map(lamdaA => P(1)(35),lamdaB => P(1)(291),lamdaOut => P(0)(35));
F136: entity F port map(lamdaA => P(1)(36),lamdaB => P(1)(292),lamdaOut => P(0)(36));
F137: entity F port map(lamdaA => P(1)(37),lamdaB => P(1)(293),lamdaOut => P(0)(37));
F138: entity F port map(lamdaA => P(1)(38),lamdaB => P(1)(294),lamdaOut => P(0)(38));
F139: entity F port map(lamdaA => P(1)(39),lamdaB => P(1)(295),lamdaOut => P(0)(39));
F140: entity F port map(lamdaA => P(1)(40),lamdaB => P(1)(296),lamdaOut => P(0)(40));
F141: entity F port map(lamdaA => P(1)(41),lamdaB => P(1)(297),lamdaOut => P(0)(41));
F142: entity F port map(lamdaA => P(1)(42),lamdaB => P(1)(298),lamdaOut => P(0)(42));
F143: entity F port map(lamdaA => P(1)(43),lamdaB => P(1)(299),lamdaOut => P(0)(43));
F144: entity F port map(lamdaA => P(1)(44),lamdaB => P(1)(300),lamdaOut => P(0)(44));
F145: entity F port map(lamdaA => P(1)(45),lamdaB => P(1)(301),lamdaOut => P(0)(45));
F146: entity F port map(lamdaA => P(1)(46),lamdaB => P(1)(302),lamdaOut => P(0)(46));
F147: entity F port map(lamdaA => P(1)(47),lamdaB => P(1)(303),lamdaOut => P(0)(47));
F148: entity F port map(lamdaA => P(1)(48),lamdaB => P(1)(304),lamdaOut => P(0)(48));
F149: entity F port map(lamdaA => P(1)(49),lamdaB => P(1)(305),lamdaOut => P(0)(49));
F150: entity F port map(lamdaA => P(1)(50),lamdaB => P(1)(306),lamdaOut => P(0)(50));
F151: entity F port map(lamdaA => P(1)(51),lamdaB => P(1)(307),lamdaOut => P(0)(51));
F152: entity F port map(lamdaA => P(1)(52),lamdaB => P(1)(308),lamdaOut => P(0)(52));
F153: entity F port map(lamdaA => P(1)(53),lamdaB => P(1)(309),lamdaOut => P(0)(53));
F154: entity F port map(lamdaA => P(1)(54),lamdaB => P(1)(310),lamdaOut => P(0)(54));
F155: entity F port map(lamdaA => P(1)(55),lamdaB => P(1)(311),lamdaOut => P(0)(55));
F156: entity F port map(lamdaA => P(1)(56),lamdaB => P(1)(312),lamdaOut => P(0)(56));
F157: entity F port map(lamdaA => P(1)(57),lamdaB => P(1)(313),lamdaOut => P(0)(57));
F158: entity F port map(lamdaA => P(1)(58),lamdaB => P(1)(314),lamdaOut => P(0)(58));
F159: entity F port map(lamdaA => P(1)(59),lamdaB => P(1)(315),lamdaOut => P(0)(59));
F160: entity F port map(lamdaA => P(1)(60),lamdaB => P(1)(316),lamdaOut => P(0)(60));
F161: entity F port map(lamdaA => P(1)(61),lamdaB => P(1)(317),lamdaOut => P(0)(61));
F162: entity F port map(lamdaA => P(1)(62),lamdaB => P(1)(318),lamdaOut => P(0)(62));
F163: entity F port map(lamdaA => P(1)(63),lamdaB => P(1)(319),lamdaOut => P(0)(63));
F164: entity F port map(lamdaA => P(1)(64),lamdaB => P(1)(320),lamdaOut => P(0)(64));
F165: entity F port map(lamdaA => P(1)(65),lamdaB => P(1)(321),lamdaOut => P(0)(65));
F166: entity F port map(lamdaA => P(1)(66),lamdaB => P(1)(322),lamdaOut => P(0)(66));
F167: entity F port map(lamdaA => P(1)(67),lamdaB => P(1)(323),lamdaOut => P(0)(67));
F168: entity F port map(lamdaA => P(1)(68),lamdaB => P(1)(324),lamdaOut => P(0)(68));
F169: entity F port map(lamdaA => P(1)(69),lamdaB => P(1)(325),lamdaOut => P(0)(69));
F170: entity F port map(lamdaA => P(1)(70),lamdaB => P(1)(326),lamdaOut => P(0)(70));
F171: entity F port map(lamdaA => P(1)(71),lamdaB => P(1)(327),lamdaOut => P(0)(71));
F172: entity F port map(lamdaA => P(1)(72),lamdaB => P(1)(328),lamdaOut => P(0)(72));
F173: entity F port map(lamdaA => P(1)(73),lamdaB => P(1)(329),lamdaOut => P(0)(73));
F174: entity F port map(lamdaA => P(1)(74),lamdaB => P(1)(330),lamdaOut => P(0)(74));
F175: entity F port map(lamdaA => P(1)(75),lamdaB => P(1)(331),lamdaOut => P(0)(75));
F176: entity F port map(lamdaA => P(1)(76),lamdaB => P(1)(332),lamdaOut => P(0)(76));
F177: entity F port map(lamdaA => P(1)(77),lamdaB => P(1)(333),lamdaOut => P(0)(77));
F178: entity F port map(lamdaA => P(1)(78),lamdaB => P(1)(334),lamdaOut => P(0)(78));
F179: entity F port map(lamdaA => P(1)(79),lamdaB => P(1)(335),lamdaOut => P(0)(79));
F180: entity F port map(lamdaA => P(1)(80),lamdaB => P(1)(336),lamdaOut => P(0)(80));
F181: entity F port map(lamdaA => P(1)(81),lamdaB => P(1)(337),lamdaOut => P(0)(81));
F182: entity F port map(lamdaA => P(1)(82),lamdaB => P(1)(338),lamdaOut => P(0)(82));
F183: entity F port map(lamdaA => P(1)(83),lamdaB => P(1)(339),lamdaOut => P(0)(83));
F184: entity F port map(lamdaA => P(1)(84),lamdaB => P(1)(340),lamdaOut => P(0)(84));
F185: entity F port map(lamdaA => P(1)(85),lamdaB => P(1)(341),lamdaOut => P(0)(85));
F186: entity F port map(lamdaA => P(1)(86),lamdaB => P(1)(342),lamdaOut => P(0)(86));
F187: entity F port map(lamdaA => P(1)(87),lamdaB => P(1)(343),lamdaOut => P(0)(87));
F188: entity F port map(lamdaA => P(1)(88),lamdaB => P(1)(344),lamdaOut => P(0)(88));
F189: entity F port map(lamdaA => P(1)(89),lamdaB => P(1)(345),lamdaOut => P(0)(89));
F190: entity F port map(lamdaA => P(1)(90),lamdaB => P(1)(346),lamdaOut => P(0)(90));
F191: entity F port map(lamdaA => P(1)(91),lamdaB => P(1)(347),lamdaOut => P(0)(91));
F192: entity F port map(lamdaA => P(1)(92),lamdaB => P(1)(348),lamdaOut => P(0)(92));
F193: entity F port map(lamdaA => P(1)(93),lamdaB => P(1)(349),lamdaOut => P(0)(93));
F194: entity F port map(lamdaA => P(1)(94),lamdaB => P(1)(350),lamdaOut => P(0)(94));
F195: entity F port map(lamdaA => P(1)(95),lamdaB => P(1)(351),lamdaOut => P(0)(95));
F196: entity F port map(lamdaA => P(1)(96),lamdaB => P(1)(352),lamdaOut => P(0)(96));
F197: entity F port map(lamdaA => P(1)(97),lamdaB => P(1)(353),lamdaOut => P(0)(97));
F198: entity F port map(lamdaA => P(1)(98),lamdaB => P(1)(354),lamdaOut => P(0)(98));
F199: entity F port map(lamdaA => P(1)(99),lamdaB => P(1)(355),lamdaOut => P(0)(99));
F1100: entity F port map(lamdaA => P(1)(100),lamdaB => P(1)(356),lamdaOut => P(0)(100));
F1101: entity F port map(lamdaA => P(1)(101),lamdaB => P(1)(357),lamdaOut => P(0)(101));
F1102: entity F port map(lamdaA => P(1)(102),lamdaB => P(1)(358),lamdaOut => P(0)(102));
F1103: entity F port map(lamdaA => P(1)(103),lamdaB => P(1)(359),lamdaOut => P(0)(103));
F1104: entity F port map(lamdaA => P(1)(104),lamdaB => P(1)(360),lamdaOut => P(0)(104));
F1105: entity F port map(lamdaA => P(1)(105),lamdaB => P(1)(361),lamdaOut => P(0)(105));
F1106: entity F port map(lamdaA => P(1)(106),lamdaB => P(1)(362),lamdaOut => P(0)(106));
F1107: entity F port map(lamdaA => P(1)(107),lamdaB => P(1)(363),lamdaOut => P(0)(107));
F1108: entity F port map(lamdaA => P(1)(108),lamdaB => P(1)(364),lamdaOut => P(0)(108));
F1109: entity F port map(lamdaA => P(1)(109),lamdaB => P(1)(365),lamdaOut => P(0)(109));
F1110: entity F port map(lamdaA => P(1)(110),lamdaB => P(1)(366),lamdaOut => P(0)(110));
F1111: entity F port map(lamdaA => P(1)(111),lamdaB => P(1)(367),lamdaOut => P(0)(111));
F1112: entity F port map(lamdaA => P(1)(112),lamdaB => P(1)(368),lamdaOut => P(0)(112));
F1113: entity F port map(lamdaA => P(1)(113),lamdaB => P(1)(369),lamdaOut => P(0)(113));
F1114: entity F port map(lamdaA => P(1)(114),lamdaB => P(1)(370),lamdaOut => P(0)(114));
F1115: entity F port map(lamdaA => P(1)(115),lamdaB => P(1)(371),lamdaOut => P(0)(115));
F1116: entity F port map(lamdaA => P(1)(116),lamdaB => P(1)(372),lamdaOut => P(0)(116));
F1117: entity F port map(lamdaA => P(1)(117),lamdaB => P(1)(373),lamdaOut => P(0)(117));
F1118: entity F port map(lamdaA => P(1)(118),lamdaB => P(1)(374),lamdaOut => P(0)(118));
F1119: entity F port map(lamdaA => P(1)(119),lamdaB => P(1)(375),lamdaOut => P(0)(119));
F1120: entity F port map(lamdaA => P(1)(120),lamdaB => P(1)(376),lamdaOut => P(0)(120));
F1121: entity F port map(lamdaA => P(1)(121),lamdaB => P(1)(377),lamdaOut => P(0)(121));
F1122: entity F port map(lamdaA => P(1)(122),lamdaB => P(1)(378),lamdaOut => P(0)(122));
F1123: entity F port map(lamdaA => P(1)(123),lamdaB => P(1)(379),lamdaOut => P(0)(123));
F1124: entity F port map(lamdaA => P(1)(124),lamdaB => P(1)(380),lamdaOut => P(0)(124));
F1125: entity F port map(lamdaA => P(1)(125),lamdaB => P(1)(381),lamdaOut => P(0)(125));
F1126: entity F port map(lamdaA => P(1)(126),lamdaB => P(1)(382),lamdaOut => P(0)(126));
F1127: entity F port map(lamdaA => P(1)(127),lamdaB => P(1)(383),lamdaOut => P(0)(127));
F1128: entity F port map(lamdaA => P(1)(128),lamdaB => P(1)(384),lamdaOut => P(0)(128));
F1129: entity F port map(lamdaA => P(1)(129),lamdaB => P(1)(385),lamdaOut => P(0)(129));
F1130: entity F port map(lamdaA => P(1)(130),lamdaB => P(1)(386),lamdaOut => P(0)(130));
F1131: entity F port map(lamdaA => P(1)(131),lamdaB => P(1)(387),lamdaOut => P(0)(131));
F1132: entity F port map(lamdaA => P(1)(132),lamdaB => P(1)(388),lamdaOut => P(0)(132));
F1133: entity F port map(lamdaA => P(1)(133),lamdaB => P(1)(389),lamdaOut => P(0)(133));
F1134: entity F port map(lamdaA => P(1)(134),lamdaB => P(1)(390),lamdaOut => P(0)(134));
F1135: entity F port map(lamdaA => P(1)(135),lamdaB => P(1)(391),lamdaOut => P(0)(135));
F1136: entity F port map(lamdaA => P(1)(136),lamdaB => P(1)(392),lamdaOut => P(0)(136));
F1137: entity F port map(lamdaA => P(1)(137),lamdaB => P(1)(393),lamdaOut => P(0)(137));
F1138: entity F port map(lamdaA => P(1)(138),lamdaB => P(1)(394),lamdaOut => P(0)(138));
F1139: entity F port map(lamdaA => P(1)(139),lamdaB => P(1)(395),lamdaOut => P(0)(139));
F1140: entity F port map(lamdaA => P(1)(140),lamdaB => P(1)(396),lamdaOut => P(0)(140));
F1141: entity F port map(lamdaA => P(1)(141),lamdaB => P(1)(397),lamdaOut => P(0)(141));
F1142: entity F port map(lamdaA => P(1)(142),lamdaB => P(1)(398),lamdaOut => P(0)(142));
F1143: entity F port map(lamdaA => P(1)(143),lamdaB => P(1)(399),lamdaOut => P(0)(143));
F1144: entity F port map(lamdaA => P(1)(144),lamdaB => P(1)(400),lamdaOut => P(0)(144));
F1145: entity F port map(lamdaA => P(1)(145),lamdaB => P(1)(401),lamdaOut => P(0)(145));
F1146: entity F port map(lamdaA => P(1)(146),lamdaB => P(1)(402),lamdaOut => P(0)(146));
F1147: entity F port map(lamdaA => P(1)(147),lamdaB => P(1)(403),lamdaOut => P(0)(147));
F1148: entity F port map(lamdaA => P(1)(148),lamdaB => P(1)(404),lamdaOut => P(0)(148));
F1149: entity F port map(lamdaA => P(1)(149),lamdaB => P(1)(405),lamdaOut => P(0)(149));
F1150: entity F port map(lamdaA => P(1)(150),lamdaB => P(1)(406),lamdaOut => P(0)(150));
F1151: entity F port map(lamdaA => P(1)(151),lamdaB => P(1)(407),lamdaOut => P(0)(151));
F1152: entity F port map(lamdaA => P(1)(152),lamdaB => P(1)(408),lamdaOut => P(0)(152));
F1153: entity F port map(lamdaA => P(1)(153),lamdaB => P(1)(409),lamdaOut => P(0)(153));
F1154: entity F port map(lamdaA => P(1)(154),lamdaB => P(1)(410),lamdaOut => P(0)(154));
F1155: entity F port map(lamdaA => P(1)(155),lamdaB => P(1)(411),lamdaOut => P(0)(155));
F1156: entity F port map(lamdaA => P(1)(156),lamdaB => P(1)(412),lamdaOut => P(0)(156));
F1157: entity F port map(lamdaA => P(1)(157),lamdaB => P(1)(413),lamdaOut => P(0)(157));
F1158: entity F port map(lamdaA => P(1)(158),lamdaB => P(1)(414),lamdaOut => P(0)(158));
F1159: entity F port map(lamdaA => P(1)(159),lamdaB => P(1)(415),lamdaOut => P(0)(159));
F1160: entity F port map(lamdaA => P(1)(160),lamdaB => P(1)(416),lamdaOut => P(0)(160));
F1161: entity F port map(lamdaA => P(1)(161),lamdaB => P(1)(417),lamdaOut => P(0)(161));
F1162: entity F port map(lamdaA => P(1)(162),lamdaB => P(1)(418),lamdaOut => P(0)(162));
F1163: entity F port map(lamdaA => P(1)(163),lamdaB => P(1)(419),lamdaOut => P(0)(163));
F1164: entity F port map(lamdaA => P(1)(164),lamdaB => P(1)(420),lamdaOut => P(0)(164));
F1165: entity F port map(lamdaA => P(1)(165),lamdaB => P(1)(421),lamdaOut => P(0)(165));
F1166: entity F port map(lamdaA => P(1)(166),lamdaB => P(1)(422),lamdaOut => P(0)(166));
F1167: entity F port map(lamdaA => P(1)(167),lamdaB => P(1)(423),lamdaOut => P(0)(167));
F1168: entity F port map(lamdaA => P(1)(168),lamdaB => P(1)(424),lamdaOut => P(0)(168));
F1169: entity F port map(lamdaA => P(1)(169),lamdaB => P(1)(425),lamdaOut => P(0)(169));
F1170: entity F port map(lamdaA => P(1)(170),lamdaB => P(1)(426),lamdaOut => P(0)(170));
F1171: entity F port map(lamdaA => P(1)(171),lamdaB => P(1)(427),lamdaOut => P(0)(171));
F1172: entity F port map(lamdaA => P(1)(172),lamdaB => P(1)(428),lamdaOut => P(0)(172));
F1173: entity F port map(lamdaA => P(1)(173),lamdaB => P(1)(429),lamdaOut => P(0)(173));
F1174: entity F port map(lamdaA => P(1)(174),lamdaB => P(1)(430),lamdaOut => P(0)(174));
F1175: entity F port map(lamdaA => P(1)(175),lamdaB => P(1)(431),lamdaOut => P(0)(175));
F1176: entity F port map(lamdaA => P(1)(176),lamdaB => P(1)(432),lamdaOut => P(0)(176));
F1177: entity F port map(lamdaA => P(1)(177),lamdaB => P(1)(433),lamdaOut => P(0)(177));
F1178: entity F port map(lamdaA => P(1)(178),lamdaB => P(1)(434),lamdaOut => P(0)(178));
F1179: entity F port map(lamdaA => P(1)(179),lamdaB => P(1)(435),lamdaOut => P(0)(179));
F1180: entity F port map(lamdaA => P(1)(180),lamdaB => P(1)(436),lamdaOut => P(0)(180));
F1181: entity F port map(lamdaA => P(1)(181),lamdaB => P(1)(437),lamdaOut => P(0)(181));
F1182: entity F port map(lamdaA => P(1)(182),lamdaB => P(1)(438),lamdaOut => P(0)(182));
F1183: entity F port map(lamdaA => P(1)(183),lamdaB => P(1)(439),lamdaOut => P(0)(183));
F1184: entity F port map(lamdaA => P(1)(184),lamdaB => P(1)(440),lamdaOut => P(0)(184));
F1185: entity F port map(lamdaA => P(1)(185),lamdaB => P(1)(441),lamdaOut => P(0)(185));
F1186: entity F port map(lamdaA => P(1)(186),lamdaB => P(1)(442),lamdaOut => P(0)(186));
F1187: entity F port map(lamdaA => P(1)(187),lamdaB => P(1)(443),lamdaOut => P(0)(187));
F1188: entity F port map(lamdaA => P(1)(188),lamdaB => P(1)(444),lamdaOut => P(0)(188));
F1189: entity F port map(lamdaA => P(1)(189),lamdaB => P(1)(445),lamdaOut => P(0)(189));
F1190: entity F port map(lamdaA => P(1)(190),lamdaB => P(1)(446),lamdaOut => P(0)(190));
F1191: entity F port map(lamdaA => P(1)(191),lamdaB => P(1)(447),lamdaOut => P(0)(191));
F1192: entity F port map(lamdaA => P(1)(192),lamdaB => P(1)(448),lamdaOut => P(0)(192));
F1193: entity F port map(lamdaA => P(1)(193),lamdaB => P(1)(449),lamdaOut => P(0)(193));
F1194: entity F port map(lamdaA => P(1)(194),lamdaB => P(1)(450),lamdaOut => P(0)(194));
F1195: entity F port map(lamdaA => P(1)(195),lamdaB => P(1)(451),lamdaOut => P(0)(195));
F1196: entity F port map(lamdaA => P(1)(196),lamdaB => P(1)(452),lamdaOut => P(0)(196));
F1197: entity F port map(lamdaA => P(1)(197),lamdaB => P(1)(453),lamdaOut => P(0)(197));
F1198: entity F port map(lamdaA => P(1)(198),lamdaB => P(1)(454),lamdaOut => P(0)(198));
F1199: entity F port map(lamdaA => P(1)(199),lamdaB => P(1)(455),lamdaOut => P(0)(199));
F1200: entity F port map(lamdaA => P(1)(200),lamdaB => P(1)(456),lamdaOut => P(0)(200));
F1201: entity F port map(lamdaA => P(1)(201),lamdaB => P(1)(457),lamdaOut => P(0)(201));
F1202: entity F port map(lamdaA => P(1)(202),lamdaB => P(1)(458),lamdaOut => P(0)(202));
F1203: entity F port map(lamdaA => P(1)(203),lamdaB => P(1)(459),lamdaOut => P(0)(203));
F1204: entity F port map(lamdaA => P(1)(204),lamdaB => P(1)(460),lamdaOut => P(0)(204));
F1205: entity F port map(lamdaA => P(1)(205),lamdaB => P(1)(461),lamdaOut => P(0)(205));
F1206: entity F port map(lamdaA => P(1)(206),lamdaB => P(1)(462),lamdaOut => P(0)(206));
F1207: entity F port map(lamdaA => P(1)(207),lamdaB => P(1)(463),lamdaOut => P(0)(207));
F1208: entity F port map(lamdaA => P(1)(208),lamdaB => P(1)(464),lamdaOut => P(0)(208));
F1209: entity F port map(lamdaA => P(1)(209),lamdaB => P(1)(465),lamdaOut => P(0)(209));
F1210: entity F port map(lamdaA => P(1)(210),lamdaB => P(1)(466),lamdaOut => P(0)(210));
F1211: entity F port map(lamdaA => P(1)(211),lamdaB => P(1)(467),lamdaOut => P(0)(211));
F1212: entity F port map(lamdaA => P(1)(212),lamdaB => P(1)(468),lamdaOut => P(0)(212));
F1213: entity F port map(lamdaA => P(1)(213),lamdaB => P(1)(469),lamdaOut => P(0)(213));
F1214: entity F port map(lamdaA => P(1)(214),lamdaB => P(1)(470),lamdaOut => P(0)(214));
F1215: entity F port map(lamdaA => P(1)(215),lamdaB => P(1)(471),lamdaOut => P(0)(215));
F1216: entity F port map(lamdaA => P(1)(216),lamdaB => P(1)(472),lamdaOut => P(0)(216));
F1217: entity F port map(lamdaA => P(1)(217),lamdaB => P(1)(473),lamdaOut => P(0)(217));
F1218: entity F port map(lamdaA => P(1)(218),lamdaB => P(1)(474),lamdaOut => P(0)(218));
F1219: entity F port map(lamdaA => P(1)(219),lamdaB => P(1)(475),lamdaOut => P(0)(219));
F1220: entity F port map(lamdaA => P(1)(220),lamdaB => P(1)(476),lamdaOut => P(0)(220));
F1221: entity F port map(lamdaA => P(1)(221),lamdaB => P(1)(477),lamdaOut => P(0)(221));
F1222: entity F port map(lamdaA => P(1)(222),lamdaB => P(1)(478),lamdaOut => P(0)(222));
F1223: entity F port map(lamdaA => P(1)(223),lamdaB => P(1)(479),lamdaOut => P(0)(223));
F1224: entity F port map(lamdaA => P(1)(224),lamdaB => P(1)(480),lamdaOut => P(0)(224));
F1225: entity F port map(lamdaA => P(1)(225),lamdaB => P(1)(481),lamdaOut => P(0)(225));
F1226: entity F port map(lamdaA => P(1)(226),lamdaB => P(1)(482),lamdaOut => P(0)(226));
F1227: entity F port map(lamdaA => P(1)(227),lamdaB => P(1)(483),lamdaOut => P(0)(227));
F1228: entity F port map(lamdaA => P(1)(228),lamdaB => P(1)(484),lamdaOut => P(0)(228));
F1229: entity F port map(lamdaA => P(1)(229),lamdaB => P(1)(485),lamdaOut => P(0)(229));
F1230: entity F port map(lamdaA => P(1)(230),lamdaB => P(1)(486),lamdaOut => P(0)(230));
F1231: entity F port map(lamdaA => P(1)(231),lamdaB => P(1)(487),lamdaOut => P(0)(231));
F1232: entity F port map(lamdaA => P(1)(232),lamdaB => P(1)(488),lamdaOut => P(0)(232));
F1233: entity F port map(lamdaA => P(1)(233),lamdaB => P(1)(489),lamdaOut => P(0)(233));
F1234: entity F port map(lamdaA => P(1)(234),lamdaB => P(1)(490),lamdaOut => P(0)(234));
F1235: entity F port map(lamdaA => P(1)(235),lamdaB => P(1)(491),lamdaOut => P(0)(235));
F1236: entity F port map(lamdaA => P(1)(236),lamdaB => P(1)(492),lamdaOut => P(0)(236));
F1237: entity F port map(lamdaA => P(1)(237),lamdaB => P(1)(493),lamdaOut => P(0)(237));
F1238: entity F port map(lamdaA => P(1)(238),lamdaB => P(1)(494),lamdaOut => P(0)(238));
F1239: entity F port map(lamdaA => P(1)(239),lamdaB => P(1)(495),lamdaOut => P(0)(239));
F1240: entity F port map(lamdaA => P(1)(240),lamdaB => P(1)(496),lamdaOut => P(0)(240));
F1241: entity F port map(lamdaA => P(1)(241),lamdaB => P(1)(497),lamdaOut => P(0)(241));
F1242: entity F port map(lamdaA => P(1)(242),lamdaB => P(1)(498),lamdaOut => P(0)(242));
F1243: entity F port map(lamdaA => P(1)(243),lamdaB => P(1)(499),lamdaOut => P(0)(243));
F1244: entity F port map(lamdaA => P(1)(244),lamdaB => P(1)(500),lamdaOut => P(0)(244));
F1245: entity F port map(lamdaA => P(1)(245),lamdaB => P(1)(501),lamdaOut => P(0)(245));
F1246: entity F port map(lamdaA => P(1)(246),lamdaB => P(1)(502),lamdaOut => P(0)(246));
F1247: entity F port map(lamdaA => P(1)(247),lamdaB => P(1)(503),lamdaOut => P(0)(247));
F1248: entity F port map(lamdaA => P(1)(248),lamdaB => P(1)(504),lamdaOut => P(0)(248));
F1249: entity F port map(lamdaA => P(1)(249),lamdaB => P(1)(505),lamdaOut => P(0)(249));
F1250: entity F port map(lamdaA => P(1)(250),lamdaB => P(1)(506),lamdaOut => P(0)(250));
F1251: entity F port map(lamdaA => P(1)(251),lamdaB => P(1)(507),lamdaOut => P(0)(251));
F1252: entity F port map(lamdaA => P(1)(252),lamdaB => P(1)(508),lamdaOut => P(0)(252));
F1253: entity F port map(lamdaA => P(1)(253),lamdaB => P(1)(509),lamdaOut => P(0)(253));
F1254: entity F port map(lamdaA => P(1)(254),lamdaB => P(1)(510),lamdaOut => P(0)(254));
F1255: entity F port map(lamdaA => P(1)(255),lamdaB => P(1)(511),lamdaOut => P(0)(255));
G1256: entity G port map(lamdaA => P(1)(0),lamdaB => P(1)(256),s => s(1)(0),lamdaOut => P(0)(256));
G1257: entity G port map(lamdaA => P(1)(1),lamdaB => P(1)(257),s => s(1)(1),lamdaOut => P(0)(257));
G1258: entity G port map(lamdaA => P(1)(2),lamdaB => P(1)(258),s => s(1)(2),lamdaOut => P(0)(258));
G1259: entity G port map(lamdaA => P(1)(3),lamdaB => P(1)(259),s => s(1)(3),lamdaOut => P(0)(259));
G1260: entity G port map(lamdaA => P(1)(4),lamdaB => P(1)(260),s => s(1)(4),lamdaOut => P(0)(260));
G1261: entity G port map(lamdaA => P(1)(5),lamdaB => P(1)(261),s => s(1)(5),lamdaOut => P(0)(261));
G1262: entity G port map(lamdaA => P(1)(6),lamdaB => P(1)(262),s => s(1)(6),lamdaOut => P(0)(262));
G1263: entity G port map(lamdaA => P(1)(7),lamdaB => P(1)(263),s => s(1)(7),lamdaOut => P(0)(263));
G1264: entity G port map(lamdaA => P(1)(8),lamdaB => P(1)(264),s => s(1)(8),lamdaOut => P(0)(264));
G1265: entity G port map(lamdaA => P(1)(9),lamdaB => P(1)(265),s => s(1)(9),lamdaOut => P(0)(265));
G1266: entity G port map(lamdaA => P(1)(10),lamdaB => P(1)(266),s => s(1)(10),lamdaOut => P(0)(266));
G1267: entity G port map(lamdaA => P(1)(11),lamdaB => P(1)(267),s => s(1)(11),lamdaOut => P(0)(267));
G1268: entity G port map(lamdaA => P(1)(12),lamdaB => P(1)(268),s => s(1)(12),lamdaOut => P(0)(268));
G1269: entity G port map(lamdaA => P(1)(13),lamdaB => P(1)(269),s => s(1)(13),lamdaOut => P(0)(269));
G1270: entity G port map(lamdaA => P(1)(14),lamdaB => P(1)(270),s => s(1)(14),lamdaOut => P(0)(270));
G1271: entity G port map(lamdaA => P(1)(15),lamdaB => P(1)(271),s => s(1)(15),lamdaOut => P(0)(271));
G1272: entity G port map(lamdaA => P(1)(16),lamdaB => P(1)(272),s => s(1)(16),lamdaOut => P(0)(272));
G1273: entity G port map(lamdaA => P(1)(17),lamdaB => P(1)(273),s => s(1)(17),lamdaOut => P(0)(273));
G1274: entity G port map(lamdaA => P(1)(18),lamdaB => P(1)(274),s => s(1)(18),lamdaOut => P(0)(274));
G1275: entity G port map(lamdaA => P(1)(19),lamdaB => P(1)(275),s => s(1)(19),lamdaOut => P(0)(275));
G1276: entity G port map(lamdaA => P(1)(20),lamdaB => P(1)(276),s => s(1)(20),lamdaOut => P(0)(276));
G1277: entity G port map(lamdaA => P(1)(21),lamdaB => P(1)(277),s => s(1)(21),lamdaOut => P(0)(277));
G1278: entity G port map(lamdaA => P(1)(22),lamdaB => P(1)(278),s => s(1)(22),lamdaOut => P(0)(278));
G1279: entity G port map(lamdaA => P(1)(23),lamdaB => P(1)(279),s => s(1)(23),lamdaOut => P(0)(279));
G1280: entity G port map(lamdaA => P(1)(24),lamdaB => P(1)(280),s => s(1)(24),lamdaOut => P(0)(280));
G1281: entity G port map(lamdaA => P(1)(25),lamdaB => P(1)(281),s => s(1)(25),lamdaOut => P(0)(281));
G1282: entity G port map(lamdaA => P(1)(26),lamdaB => P(1)(282),s => s(1)(26),lamdaOut => P(0)(282));
G1283: entity G port map(lamdaA => P(1)(27),lamdaB => P(1)(283),s => s(1)(27),lamdaOut => P(0)(283));
G1284: entity G port map(lamdaA => P(1)(28),lamdaB => P(1)(284),s => s(1)(28),lamdaOut => P(0)(284));
G1285: entity G port map(lamdaA => P(1)(29),lamdaB => P(1)(285),s => s(1)(29),lamdaOut => P(0)(285));
G1286: entity G port map(lamdaA => P(1)(30),lamdaB => P(1)(286),s => s(1)(30),lamdaOut => P(0)(286));
G1287: entity G port map(lamdaA => P(1)(31),lamdaB => P(1)(287),s => s(1)(31),lamdaOut => P(0)(287));
G1288: entity G port map(lamdaA => P(1)(32),lamdaB => P(1)(288),s => s(1)(32),lamdaOut => P(0)(288));
G1289: entity G port map(lamdaA => P(1)(33),lamdaB => P(1)(289),s => s(1)(33),lamdaOut => P(0)(289));
G1290: entity G port map(lamdaA => P(1)(34),lamdaB => P(1)(290),s => s(1)(34),lamdaOut => P(0)(290));
G1291: entity G port map(lamdaA => P(1)(35),lamdaB => P(1)(291),s => s(1)(35),lamdaOut => P(0)(291));
G1292: entity G port map(lamdaA => P(1)(36),lamdaB => P(1)(292),s => s(1)(36),lamdaOut => P(0)(292));
G1293: entity G port map(lamdaA => P(1)(37),lamdaB => P(1)(293),s => s(1)(37),lamdaOut => P(0)(293));
G1294: entity G port map(lamdaA => P(1)(38),lamdaB => P(1)(294),s => s(1)(38),lamdaOut => P(0)(294));
G1295: entity G port map(lamdaA => P(1)(39),lamdaB => P(1)(295),s => s(1)(39),lamdaOut => P(0)(295));
G1296: entity G port map(lamdaA => P(1)(40),lamdaB => P(1)(296),s => s(1)(40),lamdaOut => P(0)(296));
G1297: entity G port map(lamdaA => P(1)(41),lamdaB => P(1)(297),s => s(1)(41),lamdaOut => P(0)(297));
G1298: entity G port map(lamdaA => P(1)(42),lamdaB => P(1)(298),s => s(1)(42),lamdaOut => P(0)(298));
G1299: entity G port map(lamdaA => P(1)(43),lamdaB => P(1)(299),s => s(1)(43),lamdaOut => P(0)(299));
G1300: entity G port map(lamdaA => P(1)(44),lamdaB => P(1)(300),s => s(1)(44),lamdaOut => P(0)(300));
G1301: entity G port map(lamdaA => P(1)(45),lamdaB => P(1)(301),s => s(1)(45),lamdaOut => P(0)(301));
G1302: entity G port map(lamdaA => P(1)(46),lamdaB => P(1)(302),s => s(1)(46),lamdaOut => P(0)(302));
G1303: entity G port map(lamdaA => P(1)(47),lamdaB => P(1)(303),s => s(1)(47),lamdaOut => P(0)(303));
G1304: entity G port map(lamdaA => P(1)(48),lamdaB => P(1)(304),s => s(1)(48),lamdaOut => P(0)(304));
G1305: entity G port map(lamdaA => P(1)(49),lamdaB => P(1)(305),s => s(1)(49),lamdaOut => P(0)(305));
G1306: entity G port map(lamdaA => P(1)(50),lamdaB => P(1)(306),s => s(1)(50),lamdaOut => P(0)(306));
G1307: entity G port map(lamdaA => P(1)(51),lamdaB => P(1)(307),s => s(1)(51),lamdaOut => P(0)(307));
G1308: entity G port map(lamdaA => P(1)(52),lamdaB => P(1)(308),s => s(1)(52),lamdaOut => P(0)(308));
G1309: entity G port map(lamdaA => P(1)(53),lamdaB => P(1)(309),s => s(1)(53),lamdaOut => P(0)(309));
G1310: entity G port map(lamdaA => P(1)(54),lamdaB => P(1)(310),s => s(1)(54),lamdaOut => P(0)(310));
G1311: entity G port map(lamdaA => P(1)(55),lamdaB => P(1)(311),s => s(1)(55),lamdaOut => P(0)(311));
G1312: entity G port map(lamdaA => P(1)(56),lamdaB => P(1)(312),s => s(1)(56),lamdaOut => P(0)(312));
G1313: entity G port map(lamdaA => P(1)(57),lamdaB => P(1)(313),s => s(1)(57),lamdaOut => P(0)(313));
G1314: entity G port map(lamdaA => P(1)(58),lamdaB => P(1)(314),s => s(1)(58),lamdaOut => P(0)(314));
G1315: entity G port map(lamdaA => P(1)(59),lamdaB => P(1)(315),s => s(1)(59),lamdaOut => P(0)(315));
G1316: entity G port map(lamdaA => P(1)(60),lamdaB => P(1)(316),s => s(1)(60),lamdaOut => P(0)(316));
G1317: entity G port map(lamdaA => P(1)(61),lamdaB => P(1)(317),s => s(1)(61),lamdaOut => P(0)(317));
G1318: entity G port map(lamdaA => P(1)(62),lamdaB => P(1)(318),s => s(1)(62),lamdaOut => P(0)(318));
G1319: entity G port map(lamdaA => P(1)(63),lamdaB => P(1)(319),s => s(1)(63),lamdaOut => P(0)(319));
G1320: entity G port map(lamdaA => P(1)(64),lamdaB => P(1)(320),s => s(1)(64),lamdaOut => P(0)(320));
G1321: entity G port map(lamdaA => P(1)(65),lamdaB => P(1)(321),s => s(1)(65),lamdaOut => P(0)(321));
G1322: entity G port map(lamdaA => P(1)(66),lamdaB => P(1)(322),s => s(1)(66),lamdaOut => P(0)(322));
G1323: entity G port map(lamdaA => P(1)(67),lamdaB => P(1)(323),s => s(1)(67),lamdaOut => P(0)(323));
G1324: entity G port map(lamdaA => P(1)(68),lamdaB => P(1)(324),s => s(1)(68),lamdaOut => P(0)(324));
G1325: entity G port map(lamdaA => P(1)(69),lamdaB => P(1)(325),s => s(1)(69),lamdaOut => P(0)(325));
G1326: entity G port map(lamdaA => P(1)(70),lamdaB => P(1)(326),s => s(1)(70),lamdaOut => P(0)(326));
G1327: entity G port map(lamdaA => P(1)(71),lamdaB => P(1)(327),s => s(1)(71),lamdaOut => P(0)(327));
G1328: entity G port map(lamdaA => P(1)(72),lamdaB => P(1)(328),s => s(1)(72),lamdaOut => P(0)(328));
G1329: entity G port map(lamdaA => P(1)(73),lamdaB => P(1)(329),s => s(1)(73),lamdaOut => P(0)(329));
G1330: entity G port map(lamdaA => P(1)(74),lamdaB => P(1)(330),s => s(1)(74),lamdaOut => P(0)(330));
G1331: entity G port map(lamdaA => P(1)(75),lamdaB => P(1)(331),s => s(1)(75),lamdaOut => P(0)(331));
G1332: entity G port map(lamdaA => P(1)(76),lamdaB => P(1)(332),s => s(1)(76),lamdaOut => P(0)(332));
G1333: entity G port map(lamdaA => P(1)(77),lamdaB => P(1)(333),s => s(1)(77),lamdaOut => P(0)(333));
G1334: entity G port map(lamdaA => P(1)(78),lamdaB => P(1)(334),s => s(1)(78),lamdaOut => P(0)(334));
G1335: entity G port map(lamdaA => P(1)(79),lamdaB => P(1)(335),s => s(1)(79),lamdaOut => P(0)(335));
G1336: entity G port map(lamdaA => P(1)(80),lamdaB => P(1)(336),s => s(1)(80),lamdaOut => P(0)(336));
G1337: entity G port map(lamdaA => P(1)(81),lamdaB => P(1)(337),s => s(1)(81),lamdaOut => P(0)(337));
G1338: entity G port map(lamdaA => P(1)(82),lamdaB => P(1)(338),s => s(1)(82),lamdaOut => P(0)(338));
G1339: entity G port map(lamdaA => P(1)(83),lamdaB => P(1)(339),s => s(1)(83),lamdaOut => P(0)(339));
G1340: entity G port map(lamdaA => P(1)(84),lamdaB => P(1)(340),s => s(1)(84),lamdaOut => P(0)(340));
G1341: entity G port map(lamdaA => P(1)(85),lamdaB => P(1)(341),s => s(1)(85),lamdaOut => P(0)(341));
G1342: entity G port map(lamdaA => P(1)(86),lamdaB => P(1)(342),s => s(1)(86),lamdaOut => P(0)(342));
G1343: entity G port map(lamdaA => P(1)(87),lamdaB => P(1)(343),s => s(1)(87),lamdaOut => P(0)(343));
G1344: entity G port map(lamdaA => P(1)(88),lamdaB => P(1)(344),s => s(1)(88),lamdaOut => P(0)(344));
G1345: entity G port map(lamdaA => P(1)(89),lamdaB => P(1)(345),s => s(1)(89),lamdaOut => P(0)(345));
G1346: entity G port map(lamdaA => P(1)(90),lamdaB => P(1)(346),s => s(1)(90),lamdaOut => P(0)(346));
G1347: entity G port map(lamdaA => P(1)(91),lamdaB => P(1)(347),s => s(1)(91),lamdaOut => P(0)(347));
G1348: entity G port map(lamdaA => P(1)(92),lamdaB => P(1)(348),s => s(1)(92),lamdaOut => P(0)(348));
G1349: entity G port map(lamdaA => P(1)(93),lamdaB => P(1)(349),s => s(1)(93),lamdaOut => P(0)(349));
G1350: entity G port map(lamdaA => P(1)(94),lamdaB => P(1)(350),s => s(1)(94),lamdaOut => P(0)(350));
G1351: entity G port map(lamdaA => P(1)(95),lamdaB => P(1)(351),s => s(1)(95),lamdaOut => P(0)(351));
G1352: entity G port map(lamdaA => P(1)(96),lamdaB => P(1)(352),s => s(1)(96),lamdaOut => P(0)(352));
G1353: entity G port map(lamdaA => P(1)(97),lamdaB => P(1)(353),s => s(1)(97),lamdaOut => P(0)(353));
G1354: entity G port map(lamdaA => P(1)(98),lamdaB => P(1)(354),s => s(1)(98),lamdaOut => P(0)(354));
G1355: entity G port map(lamdaA => P(1)(99),lamdaB => P(1)(355),s => s(1)(99),lamdaOut => P(0)(355));
G1356: entity G port map(lamdaA => P(1)(100),lamdaB => P(1)(356),s => s(1)(100),lamdaOut => P(0)(356));
G1357: entity G port map(lamdaA => P(1)(101),lamdaB => P(1)(357),s => s(1)(101),lamdaOut => P(0)(357));
G1358: entity G port map(lamdaA => P(1)(102),lamdaB => P(1)(358),s => s(1)(102),lamdaOut => P(0)(358));
G1359: entity G port map(lamdaA => P(1)(103),lamdaB => P(1)(359),s => s(1)(103),lamdaOut => P(0)(359));
G1360: entity G port map(lamdaA => P(1)(104),lamdaB => P(1)(360),s => s(1)(104),lamdaOut => P(0)(360));
G1361: entity G port map(lamdaA => P(1)(105),lamdaB => P(1)(361),s => s(1)(105),lamdaOut => P(0)(361));
G1362: entity G port map(lamdaA => P(1)(106),lamdaB => P(1)(362),s => s(1)(106),lamdaOut => P(0)(362));
G1363: entity G port map(lamdaA => P(1)(107),lamdaB => P(1)(363),s => s(1)(107),lamdaOut => P(0)(363));
G1364: entity G port map(lamdaA => P(1)(108),lamdaB => P(1)(364),s => s(1)(108),lamdaOut => P(0)(364));
G1365: entity G port map(lamdaA => P(1)(109),lamdaB => P(1)(365),s => s(1)(109),lamdaOut => P(0)(365));
G1366: entity G port map(lamdaA => P(1)(110),lamdaB => P(1)(366),s => s(1)(110),lamdaOut => P(0)(366));
G1367: entity G port map(lamdaA => P(1)(111),lamdaB => P(1)(367),s => s(1)(111),lamdaOut => P(0)(367));
G1368: entity G port map(lamdaA => P(1)(112),lamdaB => P(1)(368),s => s(1)(112),lamdaOut => P(0)(368));
G1369: entity G port map(lamdaA => P(1)(113),lamdaB => P(1)(369),s => s(1)(113),lamdaOut => P(0)(369));
G1370: entity G port map(lamdaA => P(1)(114),lamdaB => P(1)(370),s => s(1)(114),lamdaOut => P(0)(370));
G1371: entity G port map(lamdaA => P(1)(115),lamdaB => P(1)(371),s => s(1)(115),lamdaOut => P(0)(371));
G1372: entity G port map(lamdaA => P(1)(116),lamdaB => P(1)(372),s => s(1)(116),lamdaOut => P(0)(372));
G1373: entity G port map(lamdaA => P(1)(117),lamdaB => P(1)(373),s => s(1)(117),lamdaOut => P(0)(373));
G1374: entity G port map(lamdaA => P(1)(118),lamdaB => P(1)(374),s => s(1)(118),lamdaOut => P(0)(374));
G1375: entity G port map(lamdaA => P(1)(119),lamdaB => P(1)(375),s => s(1)(119),lamdaOut => P(0)(375));
G1376: entity G port map(lamdaA => P(1)(120),lamdaB => P(1)(376),s => s(1)(120),lamdaOut => P(0)(376));
G1377: entity G port map(lamdaA => P(1)(121),lamdaB => P(1)(377),s => s(1)(121),lamdaOut => P(0)(377));
G1378: entity G port map(lamdaA => P(1)(122),lamdaB => P(1)(378),s => s(1)(122),lamdaOut => P(0)(378));
G1379: entity G port map(lamdaA => P(1)(123),lamdaB => P(1)(379),s => s(1)(123),lamdaOut => P(0)(379));
G1380: entity G port map(lamdaA => P(1)(124),lamdaB => P(1)(380),s => s(1)(124),lamdaOut => P(0)(380));
G1381: entity G port map(lamdaA => P(1)(125),lamdaB => P(1)(381),s => s(1)(125),lamdaOut => P(0)(381));
G1382: entity G port map(lamdaA => P(1)(126),lamdaB => P(1)(382),s => s(1)(126),lamdaOut => P(0)(382));
G1383: entity G port map(lamdaA => P(1)(127),lamdaB => P(1)(383),s => s(1)(127),lamdaOut => P(0)(383));
G1384: entity G port map(lamdaA => P(1)(128),lamdaB => P(1)(384),s => s(1)(128),lamdaOut => P(0)(384));
G1385: entity G port map(lamdaA => P(1)(129),lamdaB => P(1)(385),s => s(1)(129),lamdaOut => P(0)(385));
G1386: entity G port map(lamdaA => P(1)(130),lamdaB => P(1)(386),s => s(1)(130),lamdaOut => P(0)(386));
G1387: entity G port map(lamdaA => P(1)(131),lamdaB => P(1)(387),s => s(1)(131),lamdaOut => P(0)(387));
G1388: entity G port map(lamdaA => P(1)(132),lamdaB => P(1)(388),s => s(1)(132),lamdaOut => P(0)(388));
G1389: entity G port map(lamdaA => P(1)(133),lamdaB => P(1)(389),s => s(1)(133),lamdaOut => P(0)(389));
G1390: entity G port map(lamdaA => P(1)(134),lamdaB => P(1)(390),s => s(1)(134),lamdaOut => P(0)(390));
G1391: entity G port map(lamdaA => P(1)(135),lamdaB => P(1)(391),s => s(1)(135),lamdaOut => P(0)(391));
G1392: entity G port map(lamdaA => P(1)(136),lamdaB => P(1)(392),s => s(1)(136),lamdaOut => P(0)(392));
G1393: entity G port map(lamdaA => P(1)(137),lamdaB => P(1)(393),s => s(1)(137),lamdaOut => P(0)(393));
G1394: entity G port map(lamdaA => P(1)(138),lamdaB => P(1)(394),s => s(1)(138),lamdaOut => P(0)(394));
G1395: entity G port map(lamdaA => P(1)(139),lamdaB => P(1)(395),s => s(1)(139),lamdaOut => P(0)(395));
G1396: entity G port map(lamdaA => P(1)(140),lamdaB => P(1)(396),s => s(1)(140),lamdaOut => P(0)(396));
G1397: entity G port map(lamdaA => P(1)(141),lamdaB => P(1)(397),s => s(1)(141),lamdaOut => P(0)(397));
G1398: entity G port map(lamdaA => P(1)(142),lamdaB => P(1)(398),s => s(1)(142),lamdaOut => P(0)(398));
G1399: entity G port map(lamdaA => P(1)(143),lamdaB => P(1)(399),s => s(1)(143),lamdaOut => P(0)(399));
G1400: entity G port map(lamdaA => P(1)(144),lamdaB => P(1)(400),s => s(1)(144),lamdaOut => P(0)(400));
G1401: entity G port map(lamdaA => P(1)(145),lamdaB => P(1)(401),s => s(1)(145),lamdaOut => P(0)(401));
G1402: entity G port map(lamdaA => P(1)(146),lamdaB => P(1)(402),s => s(1)(146),lamdaOut => P(0)(402));
G1403: entity G port map(lamdaA => P(1)(147),lamdaB => P(1)(403),s => s(1)(147),lamdaOut => P(0)(403));
G1404: entity G port map(lamdaA => P(1)(148),lamdaB => P(1)(404),s => s(1)(148),lamdaOut => P(0)(404));
G1405: entity G port map(lamdaA => P(1)(149),lamdaB => P(1)(405),s => s(1)(149),lamdaOut => P(0)(405));
G1406: entity G port map(lamdaA => P(1)(150),lamdaB => P(1)(406),s => s(1)(150),lamdaOut => P(0)(406));
G1407: entity G port map(lamdaA => P(1)(151),lamdaB => P(1)(407),s => s(1)(151),lamdaOut => P(0)(407));
G1408: entity G port map(lamdaA => P(1)(152),lamdaB => P(1)(408),s => s(1)(152),lamdaOut => P(0)(408));
G1409: entity G port map(lamdaA => P(1)(153),lamdaB => P(1)(409),s => s(1)(153),lamdaOut => P(0)(409));
G1410: entity G port map(lamdaA => P(1)(154),lamdaB => P(1)(410),s => s(1)(154),lamdaOut => P(0)(410));
G1411: entity G port map(lamdaA => P(1)(155),lamdaB => P(1)(411),s => s(1)(155),lamdaOut => P(0)(411));
G1412: entity G port map(lamdaA => P(1)(156),lamdaB => P(1)(412),s => s(1)(156),lamdaOut => P(0)(412));
G1413: entity G port map(lamdaA => P(1)(157),lamdaB => P(1)(413),s => s(1)(157),lamdaOut => P(0)(413));
G1414: entity G port map(lamdaA => P(1)(158),lamdaB => P(1)(414),s => s(1)(158),lamdaOut => P(0)(414));
G1415: entity G port map(lamdaA => P(1)(159),lamdaB => P(1)(415),s => s(1)(159),lamdaOut => P(0)(415));
G1416: entity G port map(lamdaA => P(1)(160),lamdaB => P(1)(416),s => s(1)(160),lamdaOut => P(0)(416));
G1417: entity G port map(lamdaA => P(1)(161),lamdaB => P(1)(417),s => s(1)(161),lamdaOut => P(0)(417));
G1418: entity G port map(lamdaA => P(1)(162),lamdaB => P(1)(418),s => s(1)(162),lamdaOut => P(0)(418));
G1419: entity G port map(lamdaA => P(1)(163),lamdaB => P(1)(419),s => s(1)(163),lamdaOut => P(0)(419));
G1420: entity G port map(lamdaA => P(1)(164),lamdaB => P(1)(420),s => s(1)(164),lamdaOut => P(0)(420));
G1421: entity G port map(lamdaA => P(1)(165),lamdaB => P(1)(421),s => s(1)(165),lamdaOut => P(0)(421));
G1422: entity G port map(lamdaA => P(1)(166),lamdaB => P(1)(422),s => s(1)(166),lamdaOut => P(0)(422));
G1423: entity G port map(lamdaA => P(1)(167),lamdaB => P(1)(423),s => s(1)(167),lamdaOut => P(0)(423));
G1424: entity G port map(lamdaA => P(1)(168),lamdaB => P(1)(424),s => s(1)(168),lamdaOut => P(0)(424));
G1425: entity G port map(lamdaA => P(1)(169),lamdaB => P(1)(425),s => s(1)(169),lamdaOut => P(0)(425));
G1426: entity G port map(lamdaA => P(1)(170),lamdaB => P(1)(426),s => s(1)(170),lamdaOut => P(0)(426));
G1427: entity G port map(lamdaA => P(1)(171),lamdaB => P(1)(427),s => s(1)(171),lamdaOut => P(0)(427));
G1428: entity G port map(lamdaA => P(1)(172),lamdaB => P(1)(428),s => s(1)(172),lamdaOut => P(0)(428));
G1429: entity G port map(lamdaA => P(1)(173),lamdaB => P(1)(429),s => s(1)(173),lamdaOut => P(0)(429));
G1430: entity G port map(lamdaA => P(1)(174),lamdaB => P(1)(430),s => s(1)(174),lamdaOut => P(0)(430));
G1431: entity G port map(lamdaA => P(1)(175),lamdaB => P(1)(431),s => s(1)(175),lamdaOut => P(0)(431));
G1432: entity G port map(lamdaA => P(1)(176),lamdaB => P(1)(432),s => s(1)(176),lamdaOut => P(0)(432));
G1433: entity G port map(lamdaA => P(1)(177),lamdaB => P(1)(433),s => s(1)(177),lamdaOut => P(0)(433));
G1434: entity G port map(lamdaA => P(1)(178),lamdaB => P(1)(434),s => s(1)(178),lamdaOut => P(0)(434));
G1435: entity G port map(lamdaA => P(1)(179),lamdaB => P(1)(435),s => s(1)(179),lamdaOut => P(0)(435));
G1436: entity G port map(lamdaA => P(1)(180),lamdaB => P(1)(436),s => s(1)(180),lamdaOut => P(0)(436));
G1437: entity G port map(lamdaA => P(1)(181),lamdaB => P(1)(437),s => s(1)(181),lamdaOut => P(0)(437));
G1438: entity G port map(lamdaA => P(1)(182),lamdaB => P(1)(438),s => s(1)(182),lamdaOut => P(0)(438));
G1439: entity G port map(lamdaA => P(1)(183),lamdaB => P(1)(439),s => s(1)(183),lamdaOut => P(0)(439));
G1440: entity G port map(lamdaA => P(1)(184),lamdaB => P(1)(440),s => s(1)(184),lamdaOut => P(0)(440));
G1441: entity G port map(lamdaA => P(1)(185),lamdaB => P(1)(441),s => s(1)(185),lamdaOut => P(0)(441));
G1442: entity G port map(lamdaA => P(1)(186),lamdaB => P(1)(442),s => s(1)(186),lamdaOut => P(0)(442));
G1443: entity G port map(lamdaA => P(1)(187),lamdaB => P(1)(443),s => s(1)(187),lamdaOut => P(0)(443));
G1444: entity G port map(lamdaA => P(1)(188),lamdaB => P(1)(444),s => s(1)(188),lamdaOut => P(0)(444));
G1445: entity G port map(lamdaA => P(1)(189),lamdaB => P(1)(445),s => s(1)(189),lamdaOut => P(0)(445));
G1446: entity G port map(lamdaA => P(1)(190),lamdaB => P(1)(446),s => s(1)(190),lamdaOut => P(0)(446));
G1447: entity G port map(lamdaA => P(1)(191),lamdaB => P(1)(447),s => s(1)(191),lamdaOut => P(0)(447));
G1448: entity G port map(lamdaA => P(1)(192),lamdaB => P(1)(448),s => s(1)(192),lamdaOut => P(0)(448));
G1449: entity G port map(lamdaA => P(1)(193),lamdaB => P(1)(449),s => s(1)(193),lamdaOut => P(0)(449));
G1450: entity G port map(lamdaA => P(1)(194),lamdaB => P(1)(450),s => s(1)(194),lamdaOut => P(0)(450));
G1451: entity G port map(lamdaA => P(1)(195),lamdaB => P(1)(451),s => s(1)(195),lamdaOut => P(0)(451));
G1452: entity G port map(lamdaA => P(1)(196),lamdaB => P(1)(452),s => s(1)(196),lamdaOut => P(0)(452));
G1453: entity G port map(lamdaA => P(1)(197),lamdaB => P(1)(453),s => s(1)(197),lamdaOut => P(0)(453));
G1454: entity G port map(lamdaA => P(1)(198),lamdaB => P(1)(454),s => s(1)(198),lamdaOut => P(0)(454));
G1455: entity G port map(lamdaA => P(1)(199),lamdaB => P(1)(455),s => s(1)(199),lamdaOut => P(0)(455));
G1456: entity G port map(lamdaA => P(1)(200),lamdaB => P(1)(456),s => s(1)(200),lamdaOut => P(0)(456));
G1457: entity G port map(lamdaA => P(1)(201),lamdaB => P(1)(457),s => s(1)(201),lamdaOut => P(0)(457));
G1458: entity G port map(lamdaA => P(1)(202),lamdaB => P(1)(458),s => s(1)(202),lamdaOut => P(0)(458));
G1459: entity G port map(lamdaA => P(1)(203),lamdaB => P(1)(459),s => s(1)(203),lamdaOut => P(0)(459));
G1460: entity G port map(lamdaA => P(1)(204),lamdaB => P(1)(460),s => s(1)(204),lamdaOut => P(0)(460));
G1461: entity G port map(lamdaA => P(1)(205),lamdaB => P(1)(461),s => s(1)(205),lamdaOut => P(0)(461));
G1462: entity G port map(lamdaA => P(1)(206),lamdaB => P(1)(462),s => s(1)(206),lamdaOut => P(0)(462));
G1463: entity G port map(lamdaA => P(1)(207),lamdaB => P(1)(463),s => s(1)(207),lamdaOut => P(0)(463));
G1464: entity G port map(lamdaA => P(1)(208),lamdaB => P(1)(464),s => s(1)(208),lamdaOut => P(0)(464));
G1465: entity G port map(lamdaA => P(1)(209),lamdaB => P(1)(465),s => s(1)(209),lamdaOut => P(0)(465));
G1466: entity G port map(lamdaA => P(1)(210),lamdaB => P(1)(466),s => s(1)(210),lamdaOut => P(0)(466));
G1467: entity G port map(lamdaA => P(1)(211),lamdaB => P(1)(467),s => s(1)(211),lamdaOut => P(0)(467));
G1468: entity G port map(lamdaA => P(1)(212),lamdaB => P(1)(468),s => s(1)(212),lamdaOut => P(0)(468));
G1469: entity G port map(lamdaA => P(1)(213),lamdaB => P(1)(469),s => s(1)(213),lamdaOut => P(0)(469));
G1470: entity G port map(lamdaA => P(1)(214),lamdaB => P(1)(470),s => s(1)(214),lamdaOut => P(0)(470));
G1471: entity G port map(lamdaA => P(1)(215),lamdaB => P(1)(471),s => s(1)(215),lamdaOut => P(0)(471));
G1472: entity G port map(lamdaA => P(1)(216),lamdaB => P(1)(472),s => s(1)(216),lamdaOut => P(0)(472));
G1473: entity G port map(lamdaA => P(1)(217),lamdaB => P(1)(473),s => s(1)(217),lamdaOut => P(0)(473));
G1474: entity G port map(lamdaA => P(1)(218),lamdaB => P(1)(474),s => s(1)(218),lamdaOut => P(0)(474));
G1475: entity G port map(lamdaA => P(1)(219),lamdaB => P(1)(475),s => s(1)(219),lamdaOut => P(0)(475));
G1476: entity G port map(lamdaA => P(1)(220),lamdaB => P(1)(476),s => s(1)(220),lamdaOut => P(0)(476));
G1477: entity G port map(lamdaA => P(1)(221),lamdaB => P(1)(477),s => s(1)(221),lamdaOut => P(0)(477));
G1478: entity G port map(lamdaA => P(1)(222),lamdaB => P(1)(478),s => s(1)(222),lamdaOut => P(0)(478));
G1479: entity G port map(lamdaA => P(1)(223),lamdaB => P(1)(479),s => s(1)(223),lamdaOut => P(0)(479));
G1480: entity G port map(lamdaA => P(1)(224),lamdaB => P(1)(480),s => s(1)(224),lamdaOut => P(0)(480));
G1481: entity G port map(lamdaA => P(1)(225),lamdaB => P(1)(481),s => s(1)(225),lamdaOut => P(0)(481));
G1482: entity G port map(lamdaA => P(1)(226),lamdaB => P(1)(482),s => s(1)(226),lamdaOut => P(0)(482));
G1483: entity G port map(lamdaA => P(1)(227),lamdaB => P(1)(483),s => s(1)(227),lamdaOut => P(0)(483));
G1484: entity G port map(lamdaA => P(1)(228),lamdaB => P(1)(484),s => s(1)(228),lamdaOut => P(0)(484));
G1485: entity G port map(lamdaA => P(1)(229),lamdaB => P(1)(485),s => s(1)(229),lamdaOut => P(0)(485));
G1486: entity G port map(lamdaA => P(1)(230),lamdaB => P(1)(486),s => s(1)(230),lamdaOut => P(0)(486));
G1487: entity G port map(lamdaA => P(1)(231),lamdaB => P(1)(487),s => s(1)(231),lamdaOut => P(0)(487));
G1488: entity G port map(lamdaA => P(1)(232),lamdaB => P(1)(488),s => s(1)(232),lamdaOut => P(0)(488));
G1489: entity G port map(lamdaA => P(1)(233),lamdaB => P(1)(489),s => s(1)(233),lamdaOut => P(0)(489));
G1490: entity G port map(lamdaA => P(1)(234),lamdaB => P(1)(490),s => s(1)(234),lamdaOut => P(0)(490));
G1491: entity G port map(lamdaA => P(1)(235),lamdaB => P(1)(491),s => s(1)(235),lamdaOut => P(0)(491));
G1492: entity G port map(lamdaA => P(1)(236),lamdaB => P(1)(492),s => s(1)(236),lamdaOut => P(0)(492));
G1493: entity G port map(lamdaA => P(1)(237),lamdaB => P(1)(493),s => s(1)(237),lamdaOut => P(0)(493));
G1494: entity G port map(lamdaA => P(1)(238),lamdaB => P(1)(494),s => s(1)(238),lamdaOut => P(0)(494));
G1495: entity G port map(lamdaA => P(1)(239),lamdaB => P(1)(495),s => s(1)(239),lamdaOut => P(0)(495));
G1496: entity G port map(lamdaA => P(1)(240),lamdaB => P(1)(496),s => s(1)(240),lamdaOut => P(0)(496));
G1497: entity G port map(lamdaA => P(1)(241),lamdaB => P(1)(497),s => s(1)(241),lamdaOut => P(0)(497));
G1498: entity G port map(lamdaA => P(1)(242),lamdaB => P(1)(498),s => s(1)(242),lamdaOut => P(0)(498));
G1499: entity G port map(lamdaA => P(1)(243),lamdaB => P(1)(499),s => s(1)(243),lamdaOut => P(0)(499));
G1500: entity G port map(lamdaA => P(1)(244),lamdaB => P(1)(500),s => s(1)(244),lamdaOut => P(0)(500));
G1501: entity G port map(lamdaA => P(1)(245),lamdaB => P(1)(501),s => s(1)(245),lamdaOut => P(0)(501));
G1502: entity G port map(lamdaA => P(1)(246),lamdaB => P(1)(502),s => s(1)(246),lamdaOut => P(0)(502));
G1503: entity G port map(lamdaA => P(1)(247),lamdaB => P(1)(503),s => s(1)(247),lamdaOut => P(0)(503));
G1504: entity G port map(lamdaA => P(1)(248),lamdaB => P(1)(504),s => s(1)(248),lamdaOut => P(0)(504));
G1505: entity G port map(lamdaA => P(1)(249),lamdaB => P(1)(505),s => s(1)(249),lamdaOut => P(0)(505));
G1506: entity G port map(lamdaA => P(1)(250),lamdaB => P(1)(506),s => s(1)(250),lamdaOut => P(0)(506));
G1507: entity G port map(lamdaA => P(1)(251),lamdaB => P(1)(507),s => s(1)(251),lamdaOut => P(0)(507));
G1508: entity G port map(lamdaA => P(1)(252),lamdaB => P(1)(508),s => s(1)(252),lamdaOut => P(0)(508));
G1509: entity G port map(lamdaA => P(1)(253),lamdaB => P(1)(509),s => s(1)(253),lamdaOut => P(0)(509));
G1510: entity G port map(lamdaA => P(1)(254),lamdaB => P(1)(510),s => s(1)(254),lamdaOut => P(0)(510));
G1511: entity G port map(lamdaA => P(1)(255),lamdaB => P(1)(511),s => s(1)(255),lamdaOut => P(0)(511));

--Output Registers
ce_outputs <= '1';

U_D_FF0: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(492)(sign_bit),
q => outputs(0));

U_D_FF1: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(476)(sign_bit),
q => outputs(1));

U_D_FF2: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(444)(sign_bit),
q => outputs(2));

U_D_FF3: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(124)(sign_bit),
q => outputs(3));

U_D_FF4: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(380)(sign_bit),
q => outputs(4));

U_D_FF5: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(252)(sign_bit),
q => outputs(5));

U_D_FF6: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(508)(sign_bit),
q => outputs(6));

U_D_FF7: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(498)(sign_bit),
q => outputs(7));

U_D_FF8: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(490)(sign_bit),
q => outputs(8));

U_D_FF9: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(346)(sign_bit),
q => outputs(9));

U_D_FF10: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(218)(sign_bit),
q => outputs(10));

U_D_FF11: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(474)(sign_bit),
q => outputs(11));

U_D_FF12: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(314)(sign_bit),
q => outputs(12));

U_D_FF13: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(186)(sign_bit),
q => outputs(13));

U_D_FF14: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(442)(sign_bit),
q => outputs(14));

U_D_FF15: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(122)(sign_bit),
q => outputs(15));

U_D_FF16: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(378)(sign_bit),
q => outputs(16));

U_D_FF17: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(250)(sign_bit),
q => outputs(17));

U_D_FF18: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(506)(sign_bit),
q => outputs(18));

U_D_FF19: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(358)(sign_bit),
q => outputs(19));

U_D_FF20: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(230)(sign_bit),
q => outputs(20));

U_D_FF21: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(486)(sign_bit),
q => outputs(21));

U_D_FF22: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(406)(sign_bit),
q => outputs(22));

U_D_FF23: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(342)(sign_bit),
q => outputs(23));

U_D_FF24: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(214)(sign_bit),
q => outputs(24));

U_D_FF25: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(470)(sign_bit),
q => outputs(25));

U_D_FF26: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(54)(sign_bit),
q => outputs(26));

U_D_FF27: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(310)(sign_bit),
q => outputs(27));

U_D_FF28: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(182)(sign_bit),
q => outputs(28));

U_D_FF29: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(438)(sign_bit),
q => outputs(29));

U_D_FF30: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(118)(sign_bit),
q => outputs(30));

U_D_FF31: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(374)(sign_bit),
q => outputs(31));

U_D_FF32: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(246)(sign_bit),
q => outputs(32));

U_D_FF33: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(502)(sign_bit),
q => outputs(33));

U_D_FF34: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(398)(sign_bit),
q => outputs(34));

U_D_FF35: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(78)(sign_bit),
q => outputs(35));

U_D_FF36: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(334)(sign_bit),
q => outputs(36));

U_D_FF37: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(206)(sign_bit),
q => outputs(37));

U_D_FF38: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(462)(sign_bit),
q => outputs(38));

U_D_FF39: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(46)(sign_bit),
q => outputs(39));

U_D_FF40: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(302)(sign_bit),
q => outputs(40));

U_D_FF41: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(174)(sign_bit),
q => outputs(41));

U_D_FF42: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(430)(sign_bit),
q => outputs(42));

U_D_FF43: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(110)(sign_bit),
q => outputs(43));

U_D_FF44: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(366)(sign_bit),
q => outputs(44));

U_D_FF45: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(238)(sign_bit),
q => outputs(45));

U_D_FF46: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(494)(sign_bit),
q => outputs(46));

U_D_FF47: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(30)(sign_bit),
q => outputs(47));

U_D_FF48: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(286)(sign_bit),
q => outputs(48));

U_D_FF49: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(158)(sign_bit),
q => outputs(49));

U_D_FF50: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(414)(sign_bit),
q => outputs(50));

U_D_FF51: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(94)(sign_bit),
q => outputs(51));

U_D_FF52: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(350)(sign_bit),
q => outputs(52));

U_D_FF53: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(222)(sign_bit),
q => outputs(53));

U_D_FF54: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(478)(sign_bit),
q => outputs(54));

U_D_FF55: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(62)(sign_bit),
q => outputs(55));

U_D_FF56: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(318)(sign_bit),
q => outputs(56));

U_D_FF57: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(190)(sign_bit),
q => outputs(57));

U_D_FF58: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(446)(sign_bit),
q => outputs(58));

U_D_FF59: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(126)(sign_bit),
q => outputs(59));

U_D_FF60: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(382)(sign_bit),
q => outputs(60));

U_D_FF61: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(254)(sign_bit),
q => outputs(61));

U_D_FF62: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(510)(sign_bit),
q => outputs(62));

U_D_FF63: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(369)(sign_bit),
q => outputs(63));

U_D_FF64: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(241)(sign_bit),
q => outputs(64));

U_D_FF65: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(497)(sign_bit),
q => outputs(65));

U_D_FF66: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(425)(sign_bit),
q => outputs(66));

U_D_FF67: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(361)(sign_bit),
q => outputs(67));

U_D_FF68: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(233)(sign_bit),
q => outputs(68));

U_D_FF69: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(489)(sign_bit),
q => outputs(69));

U_D_FF70: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(409)(sign_bit),
q => outputs(70));

U_D_FF71: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(89)(sign_bit),
q => outputs(71));

U_D_FF72: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(345)(sign_bit),
q => outputs(72));

U_D_FF73: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(217)(sign_bit),
q => outputs(73));

U_D_FF74: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(473)(sign_bit),
q => outputs(74));

U_D_FF75: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(57)(sign_bit),
q => outputs(75));

U_D_FF76: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(313)(sign_bit),
q => outputs(76));

U_D_FF77: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(185)(sign_bit),
q => outputs(77));

U_D_FF78: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(441)(sign_bit),
q => outputs(78));

U_D_FF79: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(121)(sign_bit),
q => outputs(79));

U_D_FF80: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(377)(sign_bit),
q => outputs(80));

U_D_FF81: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(249)(sign_bit),
q => outputs(81));

U_D_FF82: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(505)(sign_bit),
q => outputs(82));

U_D_FF83: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(453)(sign_bit),
q => outputs(83));

U_D_FF84: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(421)(sign_bit),
q => outputs(84));

U_D_FF85: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(101)(sign_bit),
q => outputs(85));

U_D_FF86: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(357)(sign_bit),
q => outputs(86));

U_D_FF87: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(229)(sign_bit),
q => outputs(87));

U_D_FF88: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(485)(sign_bit),
q => outputs(88));

U_D_FF89: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(277)(sign_bit),
q => outputs(89));

U_D_FF90: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(149)(sign_bit),
q => outputs(90));

U_D_FF91: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(405)(sign_bit),
q => outputs(91));

U_D_FF92: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(85)(sign_bit),
q => outputs(92));

U_D_FF93: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(341)(sign_bit),
q => outputs(93));

U_D_FF94: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(213)(sign_bit),
q => outputs(94));

U_D_FF95: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(469)(sign_bit),
q => outputs(95));

U_D_FF96: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(53)(sign_bit),
q => outputs(96));

U_D_FF97: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(309)(sign_bit),
q => outputs(97));

U_D_FF98: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(181)(sign_bit),
q => outputs(98));

U_D_FF99: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(437)(sign_bit),
q => outputs(99));

U_D_FF100: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(117)(sign_bit),
q => outputs(100));

U_D_FF101: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(373)(sign_bit),
q => outputs(101));

U_D_FF102: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(245)(sign_bit),
q => outputs(102));

U_D_FF103: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(501)(sign_bit),
q => outputs(103));

U_D_FF104: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(269)(sign_bit),
q => outputs(104));

U_D_FF105: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(141)(sign_bit),
q => outputs(105));

U_D_FF106: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(397)(sign_bit),
q => outputs(106));

U_D_FF107: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(77)(sign_bit),
q => outputs(107));

U_D_FF108: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(333)(sign_bit),
q => outputs(108));

U_D_FF109: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(205)(sign_bit),
q => outputs(109));

U_D_FF110: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(461)(sign_bit),
q => outputs(110));

U_D_FF111: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(45)(sign_bit),
q => outputs(111));

U_D_FF112: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(301)(sign_bit),
q => outputs(112));

U_D_FF113: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(173)(sign_bit),
q => outputs(113));

U_D_FF114: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(429)(sign_bit),
q => outputs(114));

U_D_FF115: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(109)(sign_bit),
q => outputs(115));

U_D_FF116: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(365)(sign_bit),
q => outputs(116));

U_D_FF117: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(237)(sign_bit),
q => outputs(117));

U_D_FF118: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(493)(sign_bit),
q => outputs(118));

U_D_FF119: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(29)(sign_bit),
q => outputs(119));

U_D_FF120: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(285)(sign_bit),
q => outputs(120));

U_D_FF121: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(157)(sign_bit),
q => outputs(121));

U_D_FF122: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(413)(sign_bit),
q => outputs(122));

U_D_FF123: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(93)(sign_bit),
q => outputs(123));

U_D_FF124: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(349)(sign_bit),
q => outputs(124));

U_D_FF125: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(221)(sign_bit),
q => outputs(125));

U_D_FF126: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(477)(sign_bit),
q => outputs(126));

U_D_FF127: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(61)(sign_bit),
q => outputs(127));

U_D_FF128: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(317)(sign_bit),
q => outputs(128));

U_D_FF129: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(189)(sign_bit),
q => outputs(129));

U_D_FF130: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(445)(sign_bit),
q => outputs(130));

U_D_FF131: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(125)(sign_bit),
q => outputs(131));

U_D_FF132: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(381)(sign_bit),
q => outputs(132));

U_D_FF133: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(253)(sign_bit),
q => outputs(133));

U_D_FF134: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(509)(sign_bit),
q => outputs(134));

U_D_FF135: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(323)(sign_bit),
q => outputs(135));

U_D_FF136: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(195)(sign_bit),
q => outputs(136));

U_D_FF137: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(451)(sign_bit),
q => outputs(137));

U_D_FF138: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(291)(sign_bit),
q => outputs(138));

U_D_FF139: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(163)(sign_bit),
q => outputs(139));

U_D_FF140: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(419)(sign_bit),
q => outputs(140));

U_D_FF141: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(99)(sign_bit),
q => outputs(141));

U_D_FF142: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(355)(sign_bit),
q => outputs(142));

U_D_FF143: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(227)(sign_bit),
q => outputs(143));

U_D_FF144: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(483)(sign_bit),
q => outputs(144));

U_D_FF145: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(275)(sign_bit),
q => outputs(145));

U_D_FF146: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(147)(sign_bit),
q => outputs(146));

U_D_FF147: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(403)(sign_bit),
q => outputs(147));

U_D_FF148: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(83)(sign_bit),
q => outputs(148));

U_D_FF149: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(339)(sign_bit),
q => outputs(149));

U_D_FF150: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(211)(sign_bit),
q => outputs(150));

U_D_FF151: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(467)(sign_bit),
q => outputs(151));

U_D_FF152: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(51)(sign_bit),
q => outputs(152));

U_D_FF153: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(307)(sign_bit),
q => outputs(153));

U_D_FF154: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(179)(sign_bit),
q => outputs(154));

U_D_FF155: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(435)(sign_bit),
q => outputs(155));

U_D_FF156: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(115)(sign_bit),
q => outputs(156));

U_D_FF157: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(371)(sign_bit),
q => outputs(157));

U_D_FF158: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(243)(sign_bit),
q => outputs(158));

U_D_FF159: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(499)(sign_bit),
q => outputs(159));

U_D_FF160: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(11)(sign_bit),
q => outputs(160));

U_D_FF161: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(267)(sign_bit),
q => outputs(161));

U_D_FF162: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(139)(sign_bit),
q => outputs(162));

U_D_FF163: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(395)(sign_bit),
q => outputs(163));

U_D_FF164: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(75)(sign_bit),
q => outputs(164));

U_D_FF165: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(331)(sign_bit),
q => outputs(165));

U_D_FF166: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(203)(sign_bit),
q => outputs(166));

U_D_FF167: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(459)(sign_bit),
q => outputs(167));

U_D_FF168: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(43)(sign_bit),
q => outputs(168));

U_D_FF169: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(299)(sign_bit),
q => outputs(169));

U_D_FF170: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(171)(sign_bit),
q => outputs(170));

U_D_FF171: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(427)(sign_bit),
q => outputs(171));

U_D_FF172: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(107)(sign_bit),
q => outputs(172));

U_D_FF173: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(363)(sign_bit),
q => outputs(173));

U_D_FF174: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(235)(sign_bit),
q => outputs(174));

U_D_FF175: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(491)(sign_bit),
q => outputs(175));

U_D_FF176: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(27)(sign_bit),
q => outputs(176));

U_D_FF177: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(283)(sign_bit),
q => outputs(177));

U_D_FF178: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(155)(sign_bit),
q => outputs(178));

U_D_FF179: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(411)(sign_bit),
q => outputs(179));

U_D_FF180: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(91)(sign_bit),
q => outputs(180));

U_D_FF181: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(347)(sign_bit),
q => outputs(181));

U_D_FF182: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(219)(sign_bit),
q => outputs(182));

U_D_FF183: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(475)(sign_bit),
q => outputs(183));

U_D_FF184: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(59)(sign_bit),
q => outputs(184));

U_D_FF185: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(315)(sign_bit),
q => outputs(185));

U_D_FF186: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(187)(sign_bit),
q => outputs(186));

U_D_FF187: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(443)(sign_bit),
q => outputs(187));

U_D_FF188: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(123)(sign_bit),
q => outputs(188));

U_D_FF189: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(379)(sign_bit),
q => outputs(189));

U_D_FF190: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(251)(sign_bit),
q => outputs(190));

U_D_FF191: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(507)(sign_bit),
q => outputs(191));

U_D_FF192: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(7)(sign_bit),
q => outputs(192));

U_D_FF193: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(263)(sign_bit),
q => outputs(193));

U_D_FF194: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(135)(sign_bit),
q => outputs(194));

U_D_FF195: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(391)(sign_bit),
q => outputs(195));

U_D_FF196: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(71)(sign_bit),
q => outputs(196));

U_D_FF197: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(327)(sign_bit),
q => outputs(197));

U_D_FF198: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(199)(sign_bit),
q => outputs(198));

U_D_FF199: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(455)(sign_bit),
q => outputs(199));

U_D_FF200: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(39)(sign_bit),
q => outputs(200));

U_D_FF201: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(295)(sign_bit),
q => outputs(201));

U_D_FF202: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(167)(sign_bit),
q => outputs(202));

U_D_FF203: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(423)(sign_bit),
q => outputs(203));

U_D_FF204: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(103)(sign_bit),
q => outputs(204));

U_D_FF205: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(359)(sign_bit),
q => outputs(205));

U_D_FF206: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(231)(sign_bit),
q => outputs(206));

U_D_FF207: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(487)(sign_bit),
q => outputs(207));

U_D_FF208: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(23)(sign_bit),
q => outputs(208));

U_D_FF209: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(279)(sign_bit),
q => outputs(209));

U_D_FF210: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(151)(sign_bit),
q => outputs(210));

U_D_FF211: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(407)(sign_bit),
q => outputs(211));

U_D_FF212: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(87)(sign_bit),
q => outputs(212));

U_D_FF213: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(343)(sign_bit),
q => outputs(213));

U_D_FF214: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(215)(sign_bit),
q => outputs(214));

U_D_FF215: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(471)(sign_bit),
q => outputs(215));

U_D_FF216: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(55)(sign_bit),
q => outputs(216));

U_D_FF217: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(311)(sign_bit),
q => outputs(217));

U_D_FF218: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(183)(sign_bit),
q => outputs(218));

U_D_FF219: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(439)(sign_bit),
q => outputs(219));

U_D_FF220: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(119)(sign_bit),
q => outputs(220));

U_D_FF221: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(375)(sign_bit),
q => outputs(221));

U_D_FF222: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(247)(sign_bit),
q => outputs(222));

U_D_FF223: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(503)(sign_bit),
q => outputs(223));

U_D_FF224: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(15)(sign_bit),
q => outputs(224));

U_D_FF225: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(271)(sign_bit),
q => outputs(225));

U_D_FF226: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(143)(sign_bit),
q => outputs(226));

U_D_FF227: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(399)(sign_bit),
q => outputs(227));

U_D_FF228: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(79)(sign_bit),
q => outputs(228));

U_D_FF229: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(335)(sign_bit),
q => outputs(229));

U_D_FF230: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(207)(sign_bit),
q => outputs(230));

U_D_FF231: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(463)(sign_bit),
q => outputs(231));

U_D_FF232: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(47)(sign_bit),
q => outputs(232));

U_D_FF233: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(303)(sign_bit),
q => outputs(233));

U_D_FF234: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(175)(sign_bit),
q => outputs(234));

U_D_FF235: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(431)(sign_bit),
q => outputs(235));

U_D_FF236: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(111)(sign_bit),
q => outputs(236));

U_D_FF237: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(367)(sign_bit),
q => outputs(237));

U_D_FF238: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(239)(sign_bit),
q => outputs(238));

U_D_FF239: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(495)(sign_bit),
q => outputs(239));

U_D_FF240: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(31)(sign_bit),
q => outputs(240));

U_D_FF241: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(287)(sign_bit),
q => outputs(241));

U_D_FF242: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(159)(sign_bit),
q => outputs(242));

U_D_FF243: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(415)(sign_bit),
q => outputs(243));

U_D_FF244: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(95)(sign_bit),
q => outputs(244));

U_D_FF245: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(351)(sign_bit),
q => outputs(245));

U_D_FF246: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(223)(sign_bit),
q => outputs(246));

U_D_FF247: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(479)(sign_bit),
q => outputs(247));

U_D_FF248: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(63)(sign_bit),
q => outputs(248));

U_D_FF249: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(319)(sign_bit),
q => outputs(249));

U_D_FF250: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(191)(sign_bit),
q => outputs(250));

U_D_FF251: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(447)(sign_bit),
q => outputs(251));

U_D_FF252: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(127)(sign_bit),
q => outputs(252));

U_D_FF253: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(383)(sign_bit),
q => outputs(253));

U_D_FF254: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(255)(sign_bit),
q => outputs(254));

U_D_FF255: entity D_FF_1bit port map(
clk => clk,
rst => rst,
ce =>ce_outputs,
d => P(0)(511)(sign_bit),
q => outputs(255));

--Partial Sums Vector
u <=P(0)(255)(sign_bit)&P(0)(383)(sign_bit)&P(0)(127)(sign_bit)&P(0)(447)(sign_bit)&P(0)(191)(sign_bit)&P(0)(319)(sign_bit)&P(0)(63)(sign_bit)&P(0)(479)(sign_bit)&P(0)(223)(sign_bit)&P(0)(351)(sign_bit)&P(0)(95)(sign_bit)&P(0)(415)(sign_bit)&P(0)(159)(sign_bit)&P(0)(287)(sign_bit)&P(0)(31)(sign_bit)&P(0)(495)(sign_bit)&P(0)(239)(sign_bit)&P(0)(367)(sign_bit)&P(0)(111)(sign_bit)&P(0)(431)(sign_bit)&P(0)(175)(sign_bit)&P(0)(303)(sign_bit)&P(0)(47)(sign_bit)&P(0)(463)(sign_bit)&P(0)(207)(sign_bit)&P(0)(335)(sign_bit)&P(0)(79)(sign_bit)&P(0)(399)(sign_bit)&P(0)(143)(sign_bit)&P(0)(271)(sign_bit)&P(0)(15)(sign_bit)&P(0)(503)(sign_bit)&P(0)(247)(sign_bit)&P(0)(375)(sign_bit)&P(0)(119)(sign_bit)&P(0)(439)(sign_bit)&P(0)(183)(sign_bit)&P(0)(311)(sign_bit)&P(0)(55)(sign_bit)&P(0)(471)(sign_bit)&P(0)(215)(sign_bit)&P(0)(343)(sign_bit)&P(0)(87)(sign_bit)&P(0)(407)(sign_bit)&P(0)(151)(sign_bit)&P(0)(279)(sign_bit)&P(0)(23)(sign_bit)&P(0)(487)(sign_bit)&P(0)(231)(sign_bit)&P(0)(359)(sign_bit)&P(0)(103)(sign_bit)&P(0)(423)(sign_bit)&P(0)(167)(sign_bit)&P(0)(295)(sign_bit)&P(0)(39)(sign_bit)&P(0)(455)(sign_bit)&P(0)(199)(sign_bit)&P(0)(327)(sign_bit)&P(0)(71)(sign_bit)&P(0)(391)(sign_bit)&P(0)(135)(sign_bit)&P(0)(263)(sign_bit)&P(0)(7)(sign_bit)&P(0)(507)(sign_bit)&P(0)(251)(sign_bit)&P(0)(379)(sign_bit)&P(0)(123)(sign_bit)&P(0)(443)(sign_bit)&P(0)(187)(sign_bit)&P(0)(315)(sign_bit)&P(0)(59)(sign_bit)&P(0)(475)(sign_bit)&P(0)(219)(sign_bit)&P(0)(347)(sign_bit)&P(0)(91)(sign_bit)&P(0)(411)(sign_bit)&P(0)(155)(sign_bit)&P(0)(283)(sign_bit)&P(0)(27)(sign_bit)&P(0)(491)(sign_bit)&P(0)(235)(sign_bit)&P(0)(363)(sign_bit)&P(0)(107)(sign_bit)&P(0)(427)(sign_bit)&P(0)(171)(sign_bit)&P(0)(299)(sign_bit)&P(0)(43)(sign_bit)&P(0)(459)(sign_bit)&P(0)(203)(sign_bit)&P(0)(331)(sign_bit)&P(0)(75)(sign_bit)&P(0)(395)(sign_bit)&P(0)(139)(sign_bit)&P(0)(267)(sign_bit)&P(0)(11)(sign_bit)&P(0)(499)(sign_bit)&P(0)(243)(sign_bit)&P(0)(371)(sign_bit)&P(0)(115)(sign_bit)&P(0)(435)(sign_bit)&P(0)(179)(sign_bit)&P(0)(307)(sign_bit)&P(0)(51)(sign_bit)&P(0)(467)(sign_bit)&P(0)(211)(sign_bit)&P(0)(339)(sign_bit)&P(0)(83)(sign_bit)&P(0)(403)(sign_bit)&P(0)(147)(sign_bit)&P(0)(275)(sign_bit)&'0'&P(0)(483)(sign_bit)&P(0)(227)(sign_bit)&P(0)(355)(sign_bit)&P(0)(99)(sign_bit)&P(0)(419)(sign_bit)&P(0)(163)(sign_bit)&P(0)(291)(sign_bit)&'0'&P(0)(451)(sign_bit)&P(0)(195)(sign_bit)&P(0)(323)(sign_bit)&'0'&'0'&'0'&'0'&'0'&P(0)(509)(sign_bit)&P(0)(253)(sign_bit)&P(0)(381)(sign_bit)&P(0)(125)(sign_bit)&P(0)(445)(sign_bit)&P(0)(189)(sign_bit)&P(0)(317)(sign_bit)&P(0)(61)(sign_bit)&P(0)(477)(sign_bit)&P(0)(221)(sign_bit)&P(0)(349)(sign_bit)&P(0)(93)(sign_bit)&P(0)(413)(sign_bit)&P(0)(157)(sign_bit)&P(0)(285)(sign_bit)&P(0)(29)(sign_bit)&P(0)(493)(sign_bit)&P(0)(237)(sign_bit)&P(0)(365)(sign_bit)&P(0)(109)(sign_bit)&P(0)(429)(sign_bit)&P(0)(173)(sign_bit)&P(0)(301)(sign_bit)&P(0)(45)(sign_bit)&P(0)(461)(sign_bit)&P(0)(205)(sign_bit)&P(0)(333)(sign_bit)&P(0)(77)(sign_bit)&P(0)(397)(sign_bit)&P(0)(141)(sign_bit)&P(0)(269)(sign_bit)&'0'&P(0)(501)(sign_bit)&P(0)(245)(sign_bit)&P(0)(373)(sign_bit)&P(0)(117)(sign_bit)&P(0)(437)(sign_bit)&P(0)(181)(sign_bit)&P(0)(309)(sign_bit)&P(0)(53)(sign_bit)&P(0)(469)(sign_bit)&P(0)(213)(sign_bit)&P(0)(341)(sign_bit)&P(0)(85)(sign_bit)&P(0)(405)(sign_bit)&P(0)(149)(sign_bit)&P(0)(277)(sign_bit)&'0'&P(0)(485)(sign_bit)&P(0)(229)(sign_bit)&P(0)(357)(sign_bit)&P(0)(101)(sign_bit)&P(0)(421)(sign_bit)&'0'&'0'&'0'&P(0)(453)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(505)(sign_bit)&P(0)(249)(sign_bit)&P(0)(377)(sign_bit)&P(0)(121)(sign_bit)&P(0)(441)(sign_bit)&P(0)(185)(sign_bit)&P(0)(313)(sign_bit)&P(0)(57)(sign_bit)&P(0)(473)(sign_bit)&P(0)(217)(sign_bit)&P(0)(345)(sign_bit)&P(0)(89)(sign_bit)&P(0)(409)(sign_bit)&'0'&'0'&'0'&P(0)(489)(sign_bit)&P(0)(233)(sign_bit)&P(0)(361)(sign_bit)&'0'&P(0)(425)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(497)(sign_bit)&P(0)(241)(sign_bit)&P(0)(369)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(510)(sign_bit)&P(0)(254)(sign_bit)&P(0)(382)(sign_bit)&P(0)(126)(sign_bit)&P(0)(446)(sign_bit)&P(0)(190)(sign_bit)&P(0)(318)(sign_bit)&P(0)(62)(sign_bit)&P(0)(478)(sign_bit)&P(0)(222)(sign_bit)&P(0)(350)(sign_bit)&P(0)(94)(sign_bit)&P(0)(414)(sign_bit)&P(0)(158)(sign_bit)&P(0)(286)(sign_bit)&P(0)(30)(sign_bit)&P(0)(494)(sign_bit)&P(0)(238)(sign_bit)&P(0)(366)(sign_bit)&P(0)(110)(sign_bit)&P(0)(430)(sign_bit)&P(0)(174)(sign_bit)&P(0)(302)(sign_bit)&P(0)(46)(sign_bit)&P(0)(462)(sign_bit)&P(0)(206)(sign_bit)&P(0)(334)(sign_bit)&P(0)(78)(sign_bit)&P(0)(398)(sign_bit)&'0'&'0'&'0'&P(0)(502)(sign_bit)&P(0)(246)(sign_bit)&P(0)(374)(sign_bit)&P(0)(118)(sign_bit)&P(0)(438)(sign_bit)&P(0)(182)(sign_bit)&P(0)(310)(sign_bit)&P(0)(54)(sign_bit)&P(0)(470)(sign_bit)&P(0)(214)(sign_bit)&P(0)(342)(sign_bit)&'0'&P(0)(406)(sign_bit)&'0'&'0'&'0'&P(0)(486)(sign_bit)&P(0)(230)(sign_bit)&P(0)(358)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(506)(sign_bit)&P(0)(250)(sign_bit)&P(0)(378)(sign_bit)&P(0)(122)(sign_bit)&P(0)(442)(sign_bit)&P(0)(186)(sign_bit)&P(0)(314)(sign_bit)&'0'&P(0)(474)(sign_bit)&P(0)(218)(sign_bit)&P(0)(346)(sign_bit)&'0'&'0'&'0'&'0'&'0'&P(0)(490)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(498)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(508)(sign_bit)&P(0)(252)(sign_bit)&P(0)(380)(sign_bit)&P(0)(124)(sign_bit)&P(0)(444)(sign_bit)&'0'&'0'&'0'&P(0)(476)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&P(0)(492)(sign_bit)&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
--Partial Sums Entity
Partials: entity work.PartialSumGenerator port map(estimated => u,
																	partial_sums => s);

end Behavioral;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std.all;

entity synt5 is
port( 
	  address1	: in signed (5 downto 0);
	  stoixeio1	: out signed (40-1 downto 0)
);
end synt5;


architecture struct of synt5 is

    type rom_type is array (35 downto 0) of signed (39 downto 0);
    constant stoixeia : rom_type :=("0000000000000001011111001010011101110000",
"0000000000000001100000100101010001011001",
"0000000000000001100010000100010000000111",
"0000000000000001100011100111101111011001",
"0000000000000001100101010000000101011001",
"0000000000000001100110111101101101101000",
"0000000000000001101000110001000100111101",
"0000000000000001101010101010101100001111",
"0000000000000001101100101011001000011001",
"0000000000000001101110110011000100011001",
"0000000000000001110001000011001111110111",
"0000000000000001110011011100100001110101",
"0000000000000001110101111111111010101111",
"0000000000000001111000101110100011000011",
"0000000000000001111011101001110001010101",
"0000000000000001111110110011001010010001",
"0000000000000010000010001100100011010001",
"0000000000000010000101111000001011010100",
"0000000000000010001001111000101010110011",
"0000000000000010001110010001001111001000",
"0000000000000010010011000101110011111011",
"0000000000000010011000011011001110100100",
"0000000000000010011110010111100010010010",
"0000000000000010100101000010011010010011",
"0000000000000010101100100101100110000100",
"0000000000000010110101001101100100001011",
"0000000000000010111111001010111000111100",
"0000000000000011001010110010100010100011",
"0000000000000011011000011111010110111110",
"0000000000000011101000100010010101011001",
"0000000000000011101111110111010111001100",
"1111111111110000011111111100010010111011",
"1111111111111111101000111110101000101101",
"1111010101100000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000");

begin

stoixeio1<=stoixeia(to_integer((unsigned(address1))));
end struct;
